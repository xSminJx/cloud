module Rx_Top(
	
)
