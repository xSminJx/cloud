module SetBody (
	i_Clk, i_Rst,
	i_Size, i_Body_x, i_Body_y,
	i_isStart,
	o_Body_x, o_Body_y
);

	input i_Clk, i_Rst;
	input [8:0] i_Size;
	input [6:0] i_Body_x
endmodule