module Snake_Game (
    i_Clk, i_Rst,
    i_Pause, i_Push,
    o_Speed_FND0, o_Speed_FND1, o_Score_FND0, o_Score_FND1, o_Score_FND2, o_Score_FND3,
    o_hsync, o_vsync, o_red, o_blue, o_green
);
    
    input i_Clk, i_Rst;
    input [3:0] i_Push;
    input i_Pause;

    output [6:0] o_Speed_FND0, o_Speed_FND1, o_Score_FND0,
                 o_Score_FND1, o_Score_FND2, o_Score_FND3;
    output [6:0] o_Hsync, o_Vsync;
    output [3:0] o_Red, o_Blue, o_Green;

    parameter XSIZE     = 48,
              YSIZE     = 64,
              MAX_SIZE  = XSIZE*YSIZE,
              LST_CLK   = 10_000, // 원래값 : 25_000_000, 시뮬레이션 위해 10_000으로 임시 변경

              IDLE      = 3'b000,
              RUN       = 3'b001,
              CHANGE    = 3'b010,
              SETBODY   = 3'b011,
              PAUSE     = 3'b100,
              STOP      = 3'b101;

    parameter DEF_SPD   = 2,
              DEF_SIZE  = 3;

    reg [24:0] c_ClkCnt, n_ClkCnt;
    reg [5:0]  c_Body_x[0:MAX_SIZE-1], n_Body_x[0:MAX_SIZE-1], // 뱀의 몸통을 저장할 배열(큐 역할)
               c_Body_y[0:MAX_SIZE-1], n_Body_y[0:MAX_SIZE-1]; 
    reg [5:0]  c_Head_x, n_Head_x,   // 뱀의 머리 위치 저장
               c_Head_y, n_Head_y;
    reg [5:0]  c_Item_x, n_Item_x,   // 아이템 위치 저장
               c_Item_y, n_Item_y;
    reg [11:0] c_Size, n_Size;       // 뱀 크기(점수랑 같은 역할)
    reg [1:0]  c_Way, n_Way,         // 뱀이 움직였던 방향
               c_Push, n_Push;       // 조이스틱 입력 저장
    reg [2:0]  c_State, n_State;
    reg [4:0]  c_Speed, n_Speed;
    reg [4:0]  c_SpdTimeCnt, n_SpdTimeCnt; // 먹이를 먹으면 일정 시간동안 속도가 빨라지는데, 그 일정시간을 저장할 레지스터

    wire [5:0] SH_o_Head_x, SH_o_Head_y;
    wire [1:0] SH_o_Way;
    wire [5:0] SB_o_Body_x[0:MAX_SIZE-1], SB_o_Body_y[0:MAX_SIZE-1];
    
    wire isLstClk = c_ClkCnt <= LST_CLK;
    wire isEat = (n_Head_x == c_Item_x && n_Head_y == c_Item_y) && c_State == CHANGE;
    wire isGameOver = (n_Head_x == 0 || n_Head_y == 0 || n_Head_x > XSIZE + 1 || n_Head_y > YSIZE); // 그리고 몸통에 박았는지도 확인(병렬처리하셈 아니면 모듈 만들던가)
    wire isSpdDw = c_SpdTimeCnt == 16;

    //사이즈값(2진수) -> FND로 변환하는거 추가해야함(스탑워치에서 했던거 써서 모듈로 따로 분리하면 될듯)

    wire [MAX_SIZE * 6-1:0] i_Body_x_flat; // 이거 몸통 배열을 벡터로 만든건데 모듈에 넣을거임
    wire [MAX_SIZE * 6-1:0] i_Body_y_flat;
    genvar i;
    generate
        for(i=0;i<MAX_SIZE;i=i+1) begin
            assign i_Body_x_flat[i*6 +:6] = c_Body_x[i];
            assign i_Body_y_flat[i*6 +:6] = c_Body_y[i];
        end
    endgenerate


    always @(posedge i_Clk or negedge i_Rst) begin
        if(!i_Rst) begin
            c_ClkCnt     = 0;
            c_Head_x     = XSIZE >> 1;
            c_Head_y     = YSIZE >> 1;
            c_Item_x     = 0;
            c_Item_y     = 0;
            c_Size       = DEF_SIZE;
            c_Way        = 0;
            c_Push       = 0;
            c_State      = IDLE;
            c_Speed      = DEF_SPD;
            c_SpdTimeCnt = 0;

            c_Body_x[0] = c_Head_x;
            c_Body_x[1] = c_Head_x;
            c_Body_x[2] = c_Head_x;
            c_Body_y[0] = c_Head_y;
            c_Body_y[1] = c_Head_y;
            c_Body_y[2] = c_Head_y;
        end else begin
            c_ClkCnt     = n_ClkCnt;
            c_Head_x     = n_Head_x;
            c_Head_y     = n_Head_y;
            c_Size       = n_Size;
            c_Way        = n_Way;
            c_Push       = n_Push;
            c_State      = n_State;
            c_Speed      = n_Speed;
            c_SpdTimeCnt = n_SpdTimeCnt;
            //무수히 많은 c_Body대입문들...
                c_Body_x[0] = n_Body_x[0];
                c_Body_y[0] = n_Body_y[0];
                c_Body_x[1] = n_Body_x[1];
                c_Body_y[1] = n_Body_y[1];
                c_Body_x[2] = n_Body_x[2];
                c_Body_y[2] = n_Body_y[2];
                c_Body_x[3] = n_Body_x[3];
                c_Body_y[3] = n_Body_y[3];
                c_Body_x[4] = n_Body_x[4];
                c_Body_y[4] = n_Body_y[4];
                c_Body_x[5] = n_Body_x[5];
                c_Body_y[5] = n_Body_y[5];
                c_Body_x[6] = n_Body_x[6];
                c_Body_y[6] = n_Body_y[6];
                c_Body_x[7] = n_Body_x[7];
                c_Body_y[7] = n_Body_y[7];
                c_Body_x[8] = n_Body_x[8];
                c_Body_y[8] = n_Body_y[8];
                c_Body_x[9] = n_Body_x[9];
                c_Body_y[9] = n_Body_y[9];
                c_Body_x[10] = n_Body_x[10];
                c_Body_y[10] = n_Body_y[10];
                c_Body_x[11] = n_Body_x[11];
                c_Body_y[11] = n_Body_y[11];
                c_Body_x[12] = n_Body_x[12];
                c_Body_y[12] = n_Body_y[12];
                c_Body_x[13] = n_Body_x[13];
                c_Body_y[13] = n_Body_y[13];
                c_Body_x[14] = n_Body_x[14];
                c_Body_y[14] = n_Body_y[14];
                c_Body_x[15] = n_Body_x[15];
                c_Body_y[15] = n_Body_y[15];
                c_Body_x[16] = n_Body_x[16];
                c_Body_y[16] = n_Body_y[16];
                c_Body_x[17] = n_Body_x[17];
                c_Body_y[17] = n_Body_y[17];
                c_Body_x[18] = n_Body_x[18];
                c_Body_y[18] = n_Body_y[18];
                c_Body_x[19] = n_Body_x[19];
                c_Body_y[19] = n_Body_y[19];
                c_Body_x[20] = n_Body_x[20];
                c_Body_y[20] = n_Body_y[20];
                c_Body_x[21] = n_Body_x[21];
                c_Body_y[21] = n_Body_y[21];
                c_Body_x[22] = n_Body_x[22];
                c_Body_y[22] = n_Body_y[22];
                c_Body_x[23] = n_Body_x[23];
                c_Body_y[23] = n_Body_y[23];
                c_Body_x[24] = n_Body_x[24];
                c_Body_y[24] = n_Body_y[24];
                c_Body_x[25] = n_Body_x[25];
                c_Body_y[25] = n_Body_y[25];
                c_Body_x[26] = n_Body_x[26];
                c_Body_y[26] = n_Body_y[26];
                c_Body_x[27] = n_Body_x[27];
                c_Body_y[27] = n_Body_y[27];
                c_Body_x[28] = n_Body_x[28];
                c_Body_y[28] = n_Body_y[28];
                c_Body_x[29] = n_Body_x[29];
                c_Body_y[29] = n_Body_y[29];
                c_Body_x[30] = n_Body_x[30];
                c_Body_y[30] = n_Body_y[30];
                c_Body_x[31] = n_Body_x[31];
                c_Body_y[31] = n_Body_y[31];
                c_Body_x[32] = n_Body_x[32];
                c_Body_y[32] = n_Body_y[32];
                c_Body_x[33] = n_Body_x[33];
                c_Body_y[33] = n_Body_y[33];
                c_Body_x[34] = n_Body_x[34];
                c_Body_y[34] = n_Body_y[34];
                c_Body_x[35] = n_Body_x[35];
                c_Body_y[35] = n_Body_y[35];
                c_Body_x[36] = n_Body_x[36];
                c_Body_y[36] = n_Body_y[36];
                c_Body_x[37] = n_Body_x[37];
                c_Body_y[37] = n_Body_y[37];
                c_Body_x[38] = n_Body_x[38];
                c_Body_y[38] = n_Body_y[38];
                c_Body_x[39] = n_Body_x[39];
                c_Body_y[39] = n_Body_y[39];
                c_Body_x[40] = n_Body_x[40];
                c_Body_y[40] = n_Body_y[40];
                c_Body_x[41] = n_Body_x[41];
                c_Body_y[41] = n_Body_y[41];
                c_Body_x[42] = n_Body_x[42];
                c_Body_y[42] = n_Body_y[42];
                c_Body_x[43] = n_Body_x[43];
                c_Body_y[43] = n_Body_y[43];
                c_Body_x[44] = n_Body_x[44];
                c_Body_y[44] = n_Body_y[44];
                c_Body_x[45] = n_Body_x[45];
                c_Body_y[45] = n_Body_y[45];
                c_Body_x[46] = n_Body_x[46];
                c_Body_y[46] = n_Body_y[46];
                c_Body_x[47] = n_Body_x[47];
                c_Body_y[47] = n_Body_y[47];
                c_Body_x[48] = n_Body_x[48];
                c_Body_y[48] = n_Body_y[48];
                c_Body_x[49] = n_Body_x[49];
                c_Body_y[49] = n_Body_y[49];
                c_Body_x[50] = n_Body_x[50];
                c_Body_y[50] = n_Body_y[50];
                c_Body_x[51] = n_Body_x[51];
                c_Body_y[51] = n_Body_y[51];
                c_Body_x[52] = n_Body_x[52];
                c_Body_y[52] = n_Body_y[52];
                c_Body_x[53] = n_Body_x[53];
                c_Body_y[53] = n_Body_y[53];
                c_Body_x[54] = n_Body_x[54];
                c_Body_y[54] = n_Body_y[54];
                c_Body_x[55] = n_Body_x[55];
                c_Body_y[55] = n_Body_y[55];
                c_Body_x[56] = n_Body_x[56];
                c_Body_y[56] = n_Body_y[56];
                c_Body_x[57] = n_Body_x[57];
                c_Body_y[57] = n_Body_y[57];
                c_Body_x[58] = n_Body_x[58];
                c_Body_y[58] = n_Body_y[58];
                c_Body_x[59] = n_Body_x[59];
                c_Body_y[59] = n_Body_y[59];
                c_Body_x[60] = n_Body_x[60];
                c_Body_y[60] = n_Body_y[60];
                c_Body_x[61] = n_Body_x[61];
                c_Body_y[61] = n_Body_y[61];
                c_Body_x[62] = n_Body_x[62];
                c_Body_y[62] = n_Body_y[62];
                c_Body_x[63] = n_Body_x[63];
                c_Body_y[63] = n_Body_y[63];
                c_Body_x[64] = n_Body_x[64];
                c_Body_y[64] = n_Body_y[64];
                c_Body_x[65] = n_Body_x[65];
                c_Body_y[65] = n_Body_y[65];
                c_Body_x[66] = n_Body_x[66];
                c_Body_y[66] = n_Body_y[66];
                c_Body_x[67] = n_Body_x[67];
                c_Body_y[67] = n_Body_y[67];
                c_Body_x[68] = n_Body_x[68];
                c_Body_y[68] = n_Body_y[68];
                c_Body_x[69] = n_Body_x[69];
                c_Body_y[69] = n_Body_y[69];
                c_Body_x[70] = n_Body_x[70];
                c_Body_y[70] = n_Body_y[70];
                c_Body_x[71] = n_Body_x[71];
                c_Body_y[71] = n_Body_y[71];
                c_Body_x[72] = n_Body_x[72];
                c_Body_y[72] = n_Body_y[72];
                c_Body_x[73] = n_Body_x[73];
                c_Body_y[73] = n_Body_y[73];
                c_Body_x[74] = n_Body_x[74];
                c_Body_y[74] = n_Body_y[74];
                c_Body_x[75] = n_Body_x[75];
                c_Body_y[75] = n_Body_y[75];
                c_Body_x[76] = n_Body_x[76];
                c_Body_y[76] = n_Body_y[76];
                c_Body_x[77] = n_Body_x[77];
                c_Body_y[77] = n_Body_y[77];
                c_Body_x[78] = n_Body_x[78];
                c_Body_y[78] = n_Body_y[78];
                c_Body_x[79] = n_Body_x[79];
                c_Body_y[79] = n_Body_y[79];
                c_Body_x[80] = n_Body_x[80];
                c_Body_y[80] = n_Body_y[80];
                c_Body_x[81] = n_Body_x[81];
                c_Body_y[81] = n_Body_y[81];
                c_Body_x[82] = n_Body_x[82];
                c_Body_y[82] = n_Body_y[82];
                c_Body_x[83] = n_Body_x[83];
                c_Body_y[83] = n_Body_y[83];
                c_Body_x[84] = n_Body_x[84];
                c_Body_y[84] = n_Body_y[84];
                c_Body_x[85] = n_Body_x[85];
                c_Body_y[85] = n_Body_y[85];
                c_Body_x[86] = n_Body_x[86];
                c_Body_y[86] = n_Body_y[86];
                c_Body_x[87] = n_Body_x[87];
                c_Body_y[87] = n_Body_y[87];
                c_Body_x[88] = n_Body_x[88];
                c_Body_y[88] = n_Body_y[88];
                c_Body_x[89] = n_Body_x[89];
                c_Body_y[89] = n_Body_y[89];
                c_Body_x[90] = n_Body_x[90];
                c_Body_y[90] = n_Body_y[90];
                c_Body_x[91] = n_Body_x[91];
                c_Body_y[91] = n_Body_y[91];
                c_Body_x[92] = n_Body_x[92];
                c_Body_y[92] = n_Body_y[92];
                c_Body_x[93] = n_Body_x[93];
                c_Body_y[93] = n_Body_y[93];
                c_Body_x[94] = n_Body_x[94];
                c_Body_y[94] = n_Body_y[94];
                c_Body_x[95] = n_Body_x[95];
                c_Body_y[95] = n_Body_y[95];
                c_Body_x[96] = n_Body_x[96];
                c_Body_y[96] = n_Body_y[96];
                c_Body_x[97] = n_Body_x[97];
                c_Body_y[97] = n_Body_y[97];
                c_Body_x[98] = n_Body_x[98];
                c_Body_y[98] = n_Body_y[98];
                c_Body_x[99] = n_Body_x[99];
                c_Body_y[99] = n_Body_y[99];
                c_Body_x[100] = n_Body_x[100];
                c_Body_y[100] = n_Body_y[100];
                c_Body_x[101] = n_Body_x[101];
                c_Body_y[101] = n_Body_y[101];
                c_Body_x[102] = n_Body_x[102];
                c_Body_y[102] = n_Body_y[102];
                c_Body_x[103] = n_Body_x[103];
                c_Body_y[103] = n_Body_y[103];
                c_Body_x[104] = n_Body_x[104];
                c_Body_y[104] = n_Body_y[104];
                c_Body_x[105] = n_Body_x[105];
                c_Body_y[105] = n_Body_y[105];
                c_Body_x[106] = n_Body_x[106];
                c_Body_y[106] = n_Body_y[106];
                c_Body_x[107] = n_Body_x[107];
                c_Body_y[107] = n_Body_y[107];
                c_Body_x[108] = n_Body_x[108];
                c_Body_y[108] = n_Body_y[108];
                c_Body_x[109] = n_Body_x[109];
                c_Body_y[109] = n_Body_y[109];
                c_Body_x[110] = n_Body_x[110];
                c_Body_y[110] = n_Body_y[110];
                c_Body_x[111] = n_Body_x[111];
                c_Body_y[111] = n_Body_y[111];
                c_Body_x[112] = n_Body_x[112];
                c_Body_y[112] = n_Body_y[112];
                c_Body_x[113] = n_Body_x[113];
                c_Body_y[113] = n_Body_y[113];
                c_Body_x[114] = n_Body_x[114];
                c_Body_y[114] = n_Body_y[114];
                c_Body_x[115] = n_Body_x[115];
                c_Body_y[115] = n_Body_y[115];
                c_Body_x[116] = n_Body_x[116];
                c_Body_y[116] = n_Body_y[116];
                c_Body_x[117] = n_Body_x[117];
                c_Body_y[117] = n_Body_y[117];
                c_Body_x[118] = n_Body_x[118];
                c_Body_y[118] = n_Body_y[118];
                c_Body_x[119] = n_Body_x[119];
                c_Body_y[119] = n_Body_y[119];
                c_Body_x[120] = n_Body_x[120];
                c_Body_y[120] = n_Body_y[120];
                c_Body_x[121] = n_Body_x[121];
                c_Body_y[121] = n_Body_y[121];
                c_Body_x[122] = n_Body_x[122];
                c_Body_y[122] = n_Body_y[122];
                c_Body_x[123] = n_Body_x[123];
                c_Body_y[123] = n_Body_y[123];
                c_Body_x[124] = n_Body_x[124];
                c_Body_y[124] = n_Body_y[124];
                c_Body_x[125] = n_Body_x[125];
                c_Body_y[125] = n_Body_y[125];
                c_Body_x[126] = n_Body_x[126];
                c_Body_y[126] = n_Body_y[126];
                c_Body_x[127] = n_Body_x[127];
                c_Body_y[127] = n_Body_y[127];
                c_Body_x[128] = n_Body_x[128];
                c_Body_y[128] = n_Body_y[128];
                c_Body_x[129] = n_Body_x[129];
                c_Body_y[129] = n_Body_y[129];
                c_Body_x[130] = n_Body_x[130];
                c_Body_y[130] = n_Body_y[130];
                c_Body_x[131] = n_Body_x[131];
                c_Body_y[131] = n_Body_y[131];
                c_Body_x[132] = n_Body_x[132];
                c_Body_y[132] = n_Body_y[132];
                c_Body_x[133] = n_Body_x[133];
                c_Body_y[133] = n_Body_y[133];
                c_Body_x[134] = n_Body_x[134];
                c_Body_y[134] = n_Body_y[134];
                c_Body_x[135] = n_Body_x[135];
                c_Body_y[135] = n_Body_y[135];
                c_Body_x[136] = n_Body_x[136];
                c_Body_y[136] = n_Body_y[136];
                c_Body_x[137] = n_Body_x[137];
                c_Body_y[137] = n_Body_y[137];
                c_Body_x[138] = n_Body_x[138];
                c_Body_y[138] = n_Body_y[138];
                c_Body_x[139] = n_Body_x[139];
                c_Body_y[139] = n_Body_y[139];
                c_Body_x[140] = n_Body_x[140];
                c_Body_y[140] = n_Body_y[140];
                c_Body_x[141] = n_Body_x[141];
                c_Body_y[141] = n_Body_y[141];
                c_Body_x[142] = n_Body_x[142];
                c_Body_y[142] = n_Body_y[142];
                c_Body_x[143] = n_Body_x[143];
                c_Body_y[143] = n_Body_y[143];
                c_Body_x[144] = n_Body_x[144];
                c_Body_y[144] = n_Body_y[144];
                c_Body_x[145] = n_Body_x[145];
                c_Body_y[145] = n_Body_y[145];
                c_Body_x[146] = n_Body_x[146];
                c_Body_y[146] = n_Body_y[146];
                c_Body_x[147] = n_Body_x[147];
                c_Body_y[147] = n_Body_y[147];
                c_Body_x[148] = n_Body_x[148];
                c_Body_y[148] = n_Body_y[148];
                c_Body_x[149] = n_Body_x[149];
                c_Body_y[149] = n_Body_y[149];
                c_Body_x[150] = n_Body_x[150];
                c_Body_y[150] = n_Body_y[150];
                c_Body_x[151] = n_Body_x[151];
                c_Body_y[151] = n_Body_y[151];
                c_Body_x[152] = n_Body_x[152];
                c_Body_y[152] = n_Body_y[152];
                c_Body_x[153] = n_Body_x[153];
                c_Body_y[153] = n_Body_y[153];
                c_Body_x[154] = n_Body_x[154];
                c_Body_y[154] = n_Body_y[154];
                c_Body_x[155] = n_Body_x[155];
                c_Body_y[155] = n_Body_y[155];
                c_Body_x[156] = n_Body_x[156];
                c_Body_y[156] = n_Body_y[156];
                c_Body_x[157] = n_Body_x[157];
                c_Body_y[157] = n_Body_y[157];
                c_Body_x[158] = n_Body_x[158];
                c_Body_y[158] = n_Body_y[158];
                c_Body_x[159] = n_Body_x[159];
                c_Body_y[159] = n_Body_y[159];
                c_Body_x[160] = n_Body_x[160];
                c_Body_y[160] = n_Body_y[160];
                c_Body_x[161] = n_Body_x[161];
                c_Body_y[161] = n_Body_y[161];
                c_Body_x[162] = n_Body_x[162];
                c_Body_y[162] = n_Body_y[162];
                c_Body_x[163] = n_Body_x[163];
                c_Body_y[163] = n_Body_y[163];
                c_Body_x[164] = n_Body_x[164];
                c_Body_y[164] = n_Body_y[164];
                c_Body_x[165] = n_Body_x[165];
                c_Body_y[165] = n_Body_y[165];
                c_Body_x[166] = n_Body_x[166];
                c_Body_y[166] = n_Body_y[166];
                c_Body_x[167] = n_Body_x[167];
                c_Body_y[167] = n_Body_y[167];
                c_Body_x[168] = n_Body_x[168];
                c_Body_y[168] = n_Body_y[168];
                c_Body_x[169] = n_Body_x[169];
                c_Body_y[169] = n_Body_y[169];
                c_Body_x[170] = n_Body_x[170];
                c_Body_y[170] = n_Body_y[170];
                c_Body_x[171] = n_Body_x[171];
                c_Body_y[171] = n_Body_y[171];
                c_Body_x[172] = n_Body_x[172];
                c_Body_y[172] = n_Body_y[172];
                c_Body_x[173] = n_Body_x[173];
                c_Body_y[173] = n_Body_y[173];
                c_Body_x[174] = n_Body_x[174];
                c_Body_y[174] = n_Body_y[174];
                c_Body_x[175] = n_Body_x[175];
                c_Body_y[175] = n_Body_y[175];
                c_Body_x[176] = n_Body_x[176];
                c_Body_y[176] = n_Body_y[176];
                c_Body_x[177] = n_Body_x[177];
                c_Body_y[177] = n_Body_y[177];
                c_Body_x[178] = n_Body_x[178];
                c_Body_y[178] = n_Body_y[178];
                c_Body_x[179] = n_Body_x[179];
                c_Body_y[179] = n_Body_y[179];
                c_Body_x[180] = n_Body_x[180];
                c_Body_y[180] = n_Body_y[180];
                c_Body_x[181] = n_Body_x[181];
                c_Body_y[181] = n_Body_y[181];
                c_Body_x[182] = n_Body_x[182];
                c_Body_y[182] = n_Body_y[182];
                c_Body_x[183] = n_Body_x[183];
                c_Body_y[183] = n_Body_y[183];
                c_Body_x[184] = n_Body_x[184];
                c_Body_y[184] = n_Body_y[184];
                c_Body_x[185] = n_Body_x[185];
                c_Body_y[185] = n_Body_y[185];
                c_Body_x[186] = n_Body_x[186];
                c_Body_y[186] = n_Body_y[186];
                c_Body_x[187] = n_Body_x[187];
                c_Body_y[187] = n_Body_y[187];
                c_Body_x[188] = n_Body_x[188];
                c_Body_y[188] = n_Body_y[188];
                c_Body_x[189] = n_Body_x[189];
                c_Body_y[189] = n_Body_y[189];
                c_Body_x[190] = n_Body_x[190];
                c_Body_y[190] = n_Body_y[190];
                c_Body_x[191] = n_Body_x[191];
                c_Body_y[191] = n_Body_y[191];
                c_Body_x[192] = n_Body_x[192];
                c_Body_y[192] = n_Body_y[192];
                c_Body_x[193] = n_Body_x[193];
                c_Body_y[193] = n_Body_y[193];
                c_Body_x[194] = n_Body_x[194];
                c_Body_y[194] = n_Body_y[194];
                c_Body_x[195] = n_Body_x[195];
                c_Body_y[195] = n_Body_y[195];
                c_Body_x[196] = n_Body_x[196];
                c_Body_y[196] = n_Body_y[196];
                c_Body_x[197] = n_Body_x[197];
                c_Body_y[197] = n_Body_y[197];
                c_Body_x[198] = n_Body_x[198];
                c_Body_y[198] = n_Body_y[198];
                c_Body_x[199] = n_Body_x[199];
                c_Body_y[199] = n_Body_y[199];
                c_Body_x[200] = n_Body_x[200];
                c_Body_y[200] = n_Body_y[200];
                c_Body_x[201] = n_Body_x[201];
                c_Body_y[201] = n_Body_y[201];
                c_Body_x[202] = n_Body_x[202];
                c_Body_y[202] = n_Body_y[202];
                c_Body_x[203] = n_Body_x[203];
                c_Body_y[203] = n_Body_y[203];
                c_Body_x[204] = n_Body_x[204];
                c_Body_y[204] = n_Body_y[204];
                c_Body_x[205] = n_Body_x[205];
                c_Body_y[205] = n_Body_y[205];
                c_Body_x[206] = n_Body_x[206];
                c_Body_y[206] = n_Body_y[206];
                c_Body_x[207] = n_Body_x[207];
                c_Body_y[207] = n_Body_y[207];
                c_Body_x[208] = n_Body_x[208];
                c_Body_y[208] = n_Body_y[208];
                c_Body_x[209] = n_Body_x[209];
                c_Body_y[209] = n_Body_y[209];
                c_Body_x[210] = n_Body_x[210];
                c_Body_y[210] = n_Body_y[210];
                c_Body_x[211] = n_Body_x[211];
                c_Body_y[211] = n_Body_y[211];
                c_Body_x[212] = n_Body_x[212];
                c_Body_y[212] = n_Body_y[212];
                c_Body_x[213] = n_Body_x[213];
                c_Body_y[213] = n_Body_y[213];
                c_Body_x[214] = n_Body_x[214];
                c_Body_y[214] = n_Body_y[214];
                c_Body_x[215] = n_Body_x[215];
                c_Body_y[215] = n_Body_y[215];
                c_Body_x[216] = n_Body_x[216];
                c_Body_y[216] = n_Body_y[216];
                c_Body_x[217] = n_Body_x[217];
                c_Body_y[217] = n_Body_y[217];
                c_Body_x[218] = n_Body_x[218];
                c_Body_y[218] = n_Body_y[218];
                c_Body_x[219] = n_Body_x[219];
                c_Body_y[219] = n_Body_y[219];
                c_Body_x[220] = n_Body_x[220];
                c_Body_y[220] = n_Body_y[220];
                c_Body_x[221] = n_Body_x[221];
                c_Body_y[221] = n_Body_y[221];
                c_Body_x[222] = n_Body_x[222];
                c_Body_y[222] = n_Body_y[222];
                c_Body_x[223] = n_Body_x[223];
                c_Body_y[223] = n_Body_y[223];
                c_Body_x[224] = n_Body_x[224];
                c_Body_y[224] = n_Body_y[224];
                c_Body_x[225] = n_Body_x[225];
                c_Body_y[225] = n_Body_y[225];
                c_Body_x[226] = n_Body_x[226];
                c_Body_y[226] = n_Body_y[226];
                c_Body_x[227] = n_Body_x[227];
                c_Body_y[227] = n_Body_y[227];
                c_Body_x[228] = n_Body_x[228];
                c_Body_y[228] = n_Body_y[228];
                c_Body_x[229] = n_Body_x[229];
                c_Body_y[229] = n_Body_y[229];
                c_Body_x[230] = n_Body_x[230];
                c_Body_y[230] = n_Body_y[230];
                c_Body_x[231] = n_Body_x[231];
                c_Body_y[231] = n_Body_y[231];
                c_Body_x[232] = n_Body_x[232];
                c_Body_y[232] = n_Body_y[232];
                c_Body_x[233] = n_Body_x[233];
                c_Body_y[233] = n_Body_y[233];
                c_Body_x[234] = n_Body_x[234];
                c_Body_y[234] = n_Body_y[234];
                c_Body_x[235] = n_Body_x[235];
                c_Body_y[235] = n_Body_y[235];
                c_Body_x[236] = n_Body_x[236];
                c_Body_y[236] = n_Body_y[236];
                c_Body_x[237] = n_Body_x[237];
                c_Body_y[237] = n_Body_y[237];
                c_Body_x[238] = n_Body_x[238];
                c_Body_y[238] = n_Body_y[238];
                c_Body_x[239] = n_Body_x[239];
                c_Body_y[239] = n_Body_y[239];
                c_Body_x[240] = n_Body_x[240];
                c_Body_y[240] = n_Body_y[240];
                c_Body_x[241] = n_Body_x[241];
                c_Body_y[241] = n_Body_y[241];
                c_Body_x[242] = n_Body_x[242];
                c_Body_y[242] = n_Body_y[242];
                c_Body_x[243] = n_Body_x[243];
                c_Body_y[243] = n_Body_y[243];
                c_Body_x[244] = n_Body_x[244];
                c_Body_y[244] = n_Body_y[244];
                c_Body_x[245] = n_Body_x[245];
                c_Body_y[245] = n_Body_y[245];
                c_Body_x[246] = n_Body_x[246];
                c_Body_y[246] = n_Body_y[246];
                c_Body_x[247] = n_Body_x[247];
                c_Body_y[247] = n_Body_y[247];
                c_Body_x[248] = n_Body_x[248];
                c_Body_y[248] = n_Body_y[248];
                c_Body_x[249] = n_Body_x[249];
                c_Body_y[249] = n_Body_y[249];
                c_Body_x[250] = n_Body_x[250];
                c_Body_y[250] = n_Body_y[250];
                c_Body_x[251] = n_Body_x[251];
                c_Body_y[251] = n_Body_y[251];
                c_Body_x[252] = n_Body_x[252];
                c_Body_y[252] = n_Body_y[252];
                c_Body_x[253] = n_Body_x[253];
                c_Body_y[253] = n_Body_y[253];
                c_Body_x[254] = n_Body_x[254];
                c_Body_y[254] = n_Body_y[254];
                c_Body_x[255] = n_Body_x[255];
                c_Body_y[255] = n_Body_y[255];
                c_Body_x[256] = n_Body_x[256];
                c_Body_y[256] = n_Body_y[256];
                c_Body_x[257] = n_Body_x[257];
                c_Body_y[257] = n_Body_y[257];
                c_Body_x[258] = n_Body_x[258];
                c_Body_y[258] = n_Body_y[258];
                c_Body_x[259] = n_Body_x[259];
                c_Body_y[259] = n_Body_y[259];
                c_Body_x[260] = n_Body_x[260];
                c_Body_y[260] = n_Body_y[260];
                c_Body_x[261] = n_Body_x[261];
                c_Body_y[261] = n_Body_y[261];
                c_Body_x[262] = n_Body_x[262];
                c_Body_y[262] = n_Body_y[262];
                c_Body_x[263] = n_Body_x[263];
                c_Body_y[263] = n_Body_y[263];
                c_Body_x[264] = n_Body_x[264];
                c_Body_y[264] = n_Body_y[264];
                c_Body_x[265] = n_Body_x[265];
                c_Body_y[265] = n_Body_y[265];
                c_Body_x[266] = n_Body_x[266];
                c_Body_y[266] = n_Body_y[266];
                c_Body_x[267] = n_Body_x[267];
                c_Body_y[267] = n_Body_y[267];
                c_Body_x[268] = n_Body_x[268];
                c_Body_y[268] = n_Body_y[268];
                c_Body_x[269] = n_Body_x[269];
                c_Body_y[269] = n_Body_y[269];
                c_Body_x[270] = n_Body_x[270];
                c_Body_y[270] = n_Body_y[270];
                c_Body_x[271] = n_Body_x[271];
                c_Body_y[271] = n_Body_y[271];
                c_Body_x[272] = n_Body_x[272];
                c_Body_y[272] = n_Body_y[272];
                c_Body_x[273] = n_Body_x[273];
                c_Body_y[273] = n_Body_y[273];
                c_Body_x[274] = n_Body_x[274];
                c_Body_y[274] = n_Body_y[274];
                c_Body_x[275] = n_Body_x[275];
                c_Body_y[275] = n_Body_y[275];
                c_Body_x[276] = n_Body_x[276];
                c_Body_y[276] = n_Body_y[276];
                c_Body_x[277] = n_Body_x[277];
                c_Body_y[277] = n_Body_y[277];
                c_Body_x[278] = n_Body_x[278];
                c_Body_y[278] = n_Body_y[278];
                c_Body_x[279] = n_Body_x[279];
                c_Body_y[279] = n_Body_y[279];
                c_Body_x[280] = n_Body_x[280];
                c_Body_y[280] = n_Body_y[280];
                c_Body_x[281] = n_Body_x[281];
                c_Body_y[281] = n_Body_y[281];
                c_Body_x[282] = n_Body_x[282];
                c_Body_y[282] = n_Body_y[282];
                c_Body_x[283] = n_Body_x[283];
                c_Body_y[283] = n_Body_y[283];
                c_Body_x[284] = n_Body_x[284];
                c_Body_y[284] = n_Body_y[284];
                c_Body_x[285] = n_Body_x[285];
                c_Body_y[285] = n_Body_y[285];
                c_Body_x[286] = n_Body_x[286];
                c_Body_y[286] = n_Body_y[286];
                c_Body_x[287] = n_Body_x[287];
                c_Body_y[287] = n_Body_y[287];
                c_Body_x[288] = n_Body_x[288];
                c_Body_y[288] = n_Body_y[288];
                c_Body_x[289] = n_Body_x[289];
                c_Body_y[289] = n_Body_y[289];
                c_Body_x[290] = n_Body_x[290];
                c_Body_y[290] = n_Body_y[290];
                c_Body_x[291] = n_Body_x[291];
                c_Body_y[291] = n_Body_y[291];
                c_Body_x[292] = n_Body_x[292];
                c_Body_y[292] = n_Body_y[292];
                c_Body_x[293] = n_Body_x[293];
                c_Body_y[293] = n_Body_y[293];
                c_Body_x[294] = n_Body_x[294];
                c_Body_y[294] = n_Body_y[294];
                c_Body_x[295] = n_Body_x[295];
                c_Body_y[295] = n_Body_y[295];
                c_Body_x[296] = n_Body_x[296];
                c_Body_y[296] = n_Body_y[296];
                c_Body_x[297] = n_Body_x[297];
                c_Body_y[297] = n_Body_y[297];
                c_Body_x[298] = n_Body_x[298];
                c_Body_y[298] = n_Body_y[298];
                c_Body_x[299] = n_Body_x[299];
                c_Body_y[299] = n_Body_y[299];
                c_Body_x[300] = n_Body_x[300];
                c_Body_y[300] = n_Body_y[300];
                c_Body_x[301] = n_Body_x[301];
                c_Body_y[301] = n_Body_y[301];
                c_Body_x[302] = n_Body_x[302];
                c_Body_y[302] = n_Body_y[302];
                c_Body_x[303] = n_Body_x[303];
                c_Body_y[303] = n_Body_y[303];
                c_Body_x[304] = n_Body_x[304];
                c_Body_y[304] = n_Body_y[304];
                c_Body_x[305] = n_Body_x[305];
                c_Body_y[305] = n_Body_y[305];
                c_Body_x[306] = n_Body_x[306];
                c_Body_y[306] = n_Body_y[306];
                c_Body_x[307] = n_Body_x[307];
                c_Body_y[307] = n_Body_y[307];
                c_Body_x[308] = n_Body_x[308];
                c_Body_y[308] = n_Body_y[308];
                c_Body_x[309] = n_Body_x[309];
                c_Body_y[309] = n_Body_y[309];
                c_Body_x[310] = n_Body_x[310];
                c_Body_y[310] = n_Body_y[310];
                c_Body_x[311] = n_Body_x[311];
                c_Body_y[311] = n_Body_y[311];
                c_Body_x[312] = n_Body_x[312];
                c_Body_y[312] = n_Body_y[312];
                c_Body_x[313] = n_Body_x[313];
                c_Body_y[313] = n_Body_y[313];
                c_Body_x[314] = n_Body_x[314];
                c_Body_y[314] = n_Body_y[314];
                c_Body_x[315] = n_Body_x[315];
                c_Body_y[315] = n_Body_y[315];
                c_Body_x[316] = n_Body_x[316];
                c_Body_y[316] = n_Body_y[316];
                c_Body_x[317] = n_Body_x[317];
                c_Body_y[317] = n_Body_y[317];
                c_Body_x[318] = n_Body_x[318];
                c_Body_y[318] = n_Body_y[318];
                c_Body_x[319] = n_Body_x[319];
                c_Body_y[319] = n_Body_y[319];
                c_Body_x[320] = n_Body_x[320];
                c_Body_y[320] = n_Body_y[320];
                c_Body_x[321] = n_Body_x[321];
                c_Body_y[321] = n_Body_y[321];
                c_Body_x[322] = n_Body_x[322];
                c_Body_y[322] = n_Body_y[322];
                c_Body_x[323] = n_Body_x[323];
                c_Body_y[323] = n_Body_y[323];
                c_Body_x[324] = n_Body_x[324];
                c_Body_y[324] = n_Body_y[324];
                c_Body_x[325] = n_Body_x[325];
                c_Body_y[325] = n_Body_y[325];
                c_Body_x[326] = n_Body_x[326];
                c_Body_y[326] = n_Body_y[326];
                c_Body_x[327] = n_Body_x[327];
                c_Body_y[327] = n_Body_y[327];
                c_Body_x[328] = n_Body_x[328];
                c_Body_y[328] = n_Body_y[328];
                c_Body_x[329] = n_Body_x[329];
                c_Body_y[329] = n_Body_y[329];
                c_Body_x[330] = n_Body_x[330];
                c_Body_y[330] = n_Body_y[330];
                c_Body_x[331] = n_Body_x[331];
                c_Body_y[331] = n_Body_y[331];
                c_Body_x[332] = n_Body_x[332];
                c_Body_y[332] = n_Body_y[332];
                c_Body_x[333] = n_Body_x[333];
                c_Body_y[333] = n_Body_y[333];
                c_Body_x[334] = n_Body_x[334];
                c_Body_y[334] = n_Body_y[334];
                c_Body_x[335] = n_Body_x[335];
                c_Body_y[335] = n_Body_y[335];
                c_Body_x[336] = n_Body_x[336];
                c_Body_y[336] = n_Body_y[336];
                c_Body_x[337] = n_Body_x[337];
                c_Body_y[337] = n_Body_y[337];
                c_Body_x[338] = n_Body_x[338];
                c_Body_y[338] = n_Body_y[338];
                c_Body_x[339] = n_Body_x[339];
                c_Body_y[339] = n_Body_y[339];
                c_Body_x[340] = n_Body_x[340];
                c_Body_y[340] = n_Body_y[340];
                c_Body_x[341] = n_Body_x[341];
                c_Body_y[341] = n_Body_y[341];
                c_Body_x[342] = n_Body_x[342];
                c_Body_y[342] = n_Body_y[342];
                c_Body_x[343] = n_Body_x[343];
                c_Body_y[343] = n_Body_y[343];
                c_Body_x[344] = n_Body_x[344];
                c_Body_y[344] = n_Body_y[344];
                c_Body_x[345] = n_Body_x[345];
                c_Body_y[345] = n_Body_y[345];
                c_Body_x[346] = n_Body_x[346];
                c_Body_y[346] = n_Body_y[346];
                c_Body_x[347] = n_Body_x[347];
                c_Body_y[347] = n_Body_y[347];
                c_Body_x[348] = n_Body_x[348];
                c_Body_y[348] = n_Body_y[348];
                c_Body_x[349] = n_Body_x[349];
                c_Body_y[349] = n_Body_y[349];
                c_Body_x[350] = n_Body_x[350];
                c_Body_y[350] = n_Body_y[350];
                c_Body_x[351] = n_Body_x[351];
                c_Body_y[351] = n_Body_y[351];
                c_Body_x[352] = n_Body_x[352];
                c_Body_y[352] = n_Body_y[352];
                c_Body_x[353] = n_Body_x[353];
                c_Body_y[353] = n_Body_y[353];
                c_Body_x[354] = n_Body_x[354];
                c_Body_y[354] = n_Body_y[354];
                c_Body_x[355] = n_Body_x[355];
                c_Body_y[355] = n_Body_y[355];
                c_Body_x[356] = n_Body_x[356];
                c_Body_y[356] = n_Body_y[356];
                c_Body_x[357] = n_Body_x[357];
                c_Body_y[357] = n_Body_y[357];
                c_Body_x[358] = n_Body_x[358];
                c_Body_y[358] = n_Body_y[358];
                c_Body_x[359] = n_Body_x[359];
                c_Body_y[359] = n_Body_y[359];
                c_Body_x[360] = n_Body_x[360];
                c_Body_y[360] = n_Body_y[360];
                c_Body_x[361] = n_Body_x[361];
                c_Body_y[361] = n_Body_y[361];
                c_Body_x[362] = n_Body_x[362];
                c_Body_y[362] = n_Body_y[362];
                c_Body_x[363] = n_Body_x[363];
                c_Body_y[363] = n_Body_y[363];
                c_Body_x[364] = n_Body_x[364];
                c_Body_y[364] = n_Body_y[364];
                c_Body_x[365] = n_Body_x[365];
                c_Body_y[365] = n_Body_y[365];
                c_Body_x[366] = n_Body_x[366];
                c_Body_y[366] = n_Body_y[366];
                c_Body_x[367] = n_Body_x[367];
                c_Body_y[367] = n_Body_y[367];
                c_Body_x[368] = n_Body_x[368];
                c_Body_y[368] = n_Body_y[368];
                c_Body_x[369] = n_Body_x[369];
                c_Body_y[369] = n_Body_y[369];
                c_Body_x[370] = n_Body_x[370];
                c_Body_y[370] = n_Body_y[370];
                c_Body_x[371] = n_Body_x[371];
                c_Body_y[371] = n_Body_y[371];
                c_Body_x[372] = n_Body_x[372];
                c_Body_y[372] = n_Body_y[372];
                c_Body_x[373] = n_Body_x[373];
                c_Body_y[373] = n_Body_y[373];
                c_Body_x[374] = n_Body_x[374];
                c_Body_y[374] = n_Body_y[374];
                c_Body_x[375] = n_Body_x[375];
                c_Body_y[375] = n_Body_y[375];
                c_Body_x[376] = n_Body_x[376];
                c_Body_y[376] = n_Body_y[376];
                c_Body_x[377] = n_Body_x[377];
                c_Body_y[377] = n_Body_y[377];
                c_Body_x[378] = n_Body_x[378];
                c_Body_y[378] = n_Body_y[378];
                c_Body_x[379] = n_Body_x[379];
                c_Body_y[379] = n_Body_y[379];
                c_Body_x[380] = n_Body_x[380];
                c_Body_y[380] = n_Body_y[380];
                c_Body_x[381] = n_Body_x[381];
                c_Body_y[381] = n_Body_y[381];
                c_Body_x[382] = n_Body_x[382];
                c_Body_y[382] = n_Body_y[382];
                c_Body_x[383] = n_Body_x[383];
                c_Body_y[383] = n_Body_y[383];
                c_Body_x[384] = n_Body_x[384];
                c_Body_y[384] = n_Body_y[384];
                c_Body_x[385] = n_Body_x[385];
                c_Body_y[385] = n_Body_y[385];
                c_Body_x[386] = n_Body_x[386];
                c_Body_y[386] = n_Body_y[386];
                c_Body_x[387] = n_Body_x[387];
                c_Body_y[387] = n_Body_y[387];
                c_Body_x[388] = n_Body_x[388];
                c_Body_y[388] = n_Body_y[388];
                c_Body_x[389] = n_Body_x[389];
                c_Body_y[389] = n_Body_y[389];
                c_Body_x[390] = n_Body_x[390];
                c_Body_y[390] = n_Body_y[390];
                c_Body_x[391] = n_Body_x[391];
                c_Body_y[391] = n_Body_y[391];
                c_Body_x[392] = n_Body_x[392];
                c_Body_y[392] = n_Body_y[392];
                c_Body_x[393] = n_Body_x[393];
                c_Body_y[393] = n_Body_y[393];
                c_Body_x[394] = n_Body_x[394];
                c_Body_y[394] = n_Body_y[394];
                c_Body_x[395] = n_Body_x[395];
                c_Body_y[395] = n_Body_y[395];
                c_Body_x[396] = n_Body_x[396];
                c_Body_y[396] = n_Body_y[396];
                c_Body_x[397] = n_Body_x[397];
                c_Body_y[397] = n_Body_y[397];
                c_Body_x[398] = n_Body_x[398];
                c_Body_y[398] = n_Body_y[398];
                c_Body_x[399] = n_Body_x[399];
                c_Body_y[399] = n_Body_y[399];
                c_Body_x[400] = n_Body_x[400];
                c_Body_y[400] = n_Body_y[400];
                c_Body_x[401] = n_Body_x[401];
                c_Body_y[401] = n_Body_y[401];
                c_Body_x[402] = n_Body_x[402];
                c_Body_y[402] = n_Body_y[402];
                c_Body_x[403] = n_Body_x[403];
                c_Body_y[403] = n_Body_y[403];
                c_Body_x[404] = n_Body_x[404];
                c_Body_y[404] = n_Body_y[404];
                c_Body_x[405] = n_Body_x[405];
                c_Body_y[405] = n_Body_y[405];
                c_Body_x[406] = n_Body_x[406];
                c_Body_y[406] = n_Body_y[406];
                c_Body_x[407] = n_Body_x[407];
                c_Body_y[407] = n_Body_y[407];
                c_Body_x[408] = n_Body_x[408];
                c_Body_y[408] = n_Body_y[408];
                c_Body_x[409] = n_Body_x[409];
                c_Body_y[409] = n_Body_y[409];
                c_Body_x[410] = n_Body_x[410];
                c_Body_y[410] = n_Body_y[410];
                c_Body_x[411] = n_Body_x[411];
                c_Body_y[411] = n_Body_y[411];
                c_Body_x[412] = n_Body_x[412];
                c_Body_y[412] = n_Body_y[412];
                c_Body_x[413] = n_Body_x[413];
                c_Body_y[413] = n_Body_y[413];
                c_Body_x[414] = n_Body_x[414];
                c_Body_y[414] = n_Body_y[414];
                c_Body_x[415] = n_Body_x[415];
                c_Body_y[415] = n_Body_y[415];
                c_Body_x[416] = n_Body_x[416];
                c_Body_y[416] = n_Body_y[416];
                c_Body_x[417] = n_Body_x[417];
                c_Body_y[417] = n_Body_y[417];
                c_Body_x[418] = n_Body_x[418];
                c_Body_y[418] = n_Body_y[418];
                c_Body_x[419] = n_Body_x[419];
                c_Body_y[419] = n_Body_y[419];
                c_Body_x[420] = n_Body_x[420];
                c_Body_y[420] = n_Body_y[420];
                c_Body_x[421] = n_Body_x[421];
                c_Body_y[421] = n_Body_y[421];
                c_Body_x[422] = n_Body_x[422];
                c_Body_y[422] = n_Body_y[422];
                c_Body_x[423] = n_Body_x[423];
                c_Body_y[423] = n_Body_y[423];
                c_Body_x[424] = n_Body_x[424];
                c_Body_y[424] = n_Body_y[424];
                c_Body_x[425] = n_Body_x[425];
                c_Body_y[425] = n_Body_y[425];
                c_Body_x[426] = n_Body_x[426];
                c_Body_y[426] = n_Body_y[426];
                c_Body_x[427] = n_Body_x[427];
                c_Body_y[427] = n_Body_y[427];
                c_Body_x[428] = n_Body_x[428];
                c_Body_y[428] = n_Body_y[428];
                c_Body_x[429] = n_Body_x[429];
                c_Body_y[429] = n_Body_y[429];
                c_Body_x[430] = n_Body_x[430];
                c_Body_y[430] = n_Body_y[430];
                c_Body_x[431] = n_Body_x[431];
                c_Body_y[431] = n_Body_y[431];
                c_Body_x[432] = n_Body_x[432];
                c_Body_y[432] = n_Body_y[432];
                c_Body_x[433] = n_Body_x[433];
                c_Body_y[433] = n_Body_y[433];
                c_Body_x[434] = n_Body_x[434];
                c_Body_y[434] = n_Body_y[434];
                c_Body_x[435] = n_Body_x[435];
                c_Body_y[435] = n_Body_y[435];
                c_Body_x[436] = n_Body_x[436];
                c_Body_y[436] = n_Body_y[436];
                c_Body_x[437] = n_Body_x[437];
                c_Body_y[437] = n_Body_y[437];
                c_Body_x[438] = n_Body_x[438];
                c_Body_y[438] = n_Body_y[438];
                c_Body_x[439] = n_Body_x[439];
                c_Body_y[439] = n_Body_y[439];
                c_Body_x[440] = n_Body_x[440];
                c_Body_y[440] = n_Body_y[440];
                c_Body_x[441] = n_Body_x[441];
                c_Body_y[441] = n_Body_y[441];
                c_Body_x[442] = n_Body_x[442];
                c_Body_y[442] = n_Body_y[442];
                c_Body_x[443] = n_Body_x[443];
                c_Body_y[443] = n_Body_y[443];
                c_Body_x[444] = n_Body_x[444];
                c_Body_y[444] = n_Body_y[444];
                c_Body_x[445] = n_Body_x[445];
                c_Body_y[445] = n_Body_y[445];
                c_Body_x[446] = n_Body_x[446];
                c_Body_y[446] = n_Body_y[446];
                c_Body_x[447] = n_Body_x[447];
                c_Body_y[447] = n_Body_y[447];
                c_Body_x[448] = n_Body_x[448];
                c_Body_y[448] = n_Body_y[448];
                c_Body_x[449] = n_Body_x[449];
                c_Body_y[449] = n_Body_y[449];
                c_Body_x[450] = n_Body_x[450];
                c_Body_y[450] = n_Body_y[450];
                c_Body_x[451] = n_Body_x[451];
                c_Body_y[451] = n_Body_y[451];
                c_Body_x[452] = n_Body_x[452];
                c_Body_y[452] = n_Body_y[452];
                c_Body_x[453] = n_Body_x[453];
                c_Body_y[453] = n_Body_y[453];
                c_Body_x[454] = n_Body_x[454];
                c_Body_y[454] = n_Body_y[454];
                c_Body_x[455] = n_Body_x[455];
                c_Body_y[455] = n_Body_y[455];
                c_Body_x[456] = n_Body_x[456];
                c_Body_y[456] = n_Body_y[456];
                c_Body_x[457] = n_Body_x[457];
                c_Body_y[457] = n_Body_y[457];
                c_Body_x[458] = n_Body_x[458];
                c_Body_y[458] = n_Body_y[458];
                c_Body_x[459] = n_Body_x[459];
                c_Body_y[459] = n_Body_y[459];
                c_Body_x[460] = n_Body_x[460];
                c_Body_y[460] = n_Body_y[460];
                c_Body_x[461] = n_Body_x[461];
                c_Body_y[461] = n_Body_y[461];
                c_Body_x[462] = n_Body_x[462];
                c_Body_y[462] = n_Body_y[462];
                c_Body_x[463] = n_Body_x[463];
                c_Body_y[463] = n_Body_y[463];
                c_Body_x[464] = n_Body_x[464];
                c_Body_y[464] = n_Body_y[464];
                c_Body_x[465] = n_Body_x[465];
                c_Body_y[465] = n_Body_y[465];
                c_Body_x[466] = n_Body_x[466];
                c_Body_y[466] = n_Body_y[466];
                c_Body_x[467] = n_Body_x[467];
                c_Body_y[467] = n_Body_y[467];
                c_Body_x[468] = n_Body_x[468];
                c_Body_y[468] = n_Body_y[468];
                c_Body_x[469] = n_Body_x[469];
                c_Body_y[469] = n_Body_y[469];
                c_Body_x[470] = n_Body_x[470];
                c_Body_y[470] = n_Body_y[470];
                c_Body_x[471] = n_Body_x[471];
                c_Body_y[471] = n_Body_y[471];
                c_Body_x[472] = n_Body_x[472];
                c_Body_y[472] = n_Body_y[472];
                c_Body_x[473] = n_Body_x[473];
                c_Body_y[473] = n_Body_y[473];
                c_Body_x[474] = n_Body_x[474];
                c_Body_y[474] = n_Body_y[474];
                c_Body_x[475] = n_Body_x[475];
                c_Body_y[475] = n_Body_y[475];
                c_Body_x[476] = n_Body_x[476];
                c_Body_y[476] = n_Body_y[476];
                c_Body_x[477] = n_Body_x[477];
                c_Body_y[477] = n_Body_y[477];
                c_Body_x[478] = n_Body_x[478];
                c_Body_y[478] = n_Body_y[478];
                c_Body_x[479] = n_Body_x[479];
                c_Body_y[479] = n_Body_y[479];
                c_Body_x[480] = n_Body_x[480];
                c_Body_y[480] = n_Body_y[480];
                c_Body_x[481] = n_Body_x[481];
                c_Body_y[481] = n_Body_y[481];
                c_Body_x[482] = n_Body_x[482];
                c_Body_y[482] = n_Body_y[482];
                c_Body_x[483] = n_Body_x[483];
                c_Body_y[483] = n_Body_y[483];
                c_Body_x[484] = n_Body_x[484];
                c_Body_y[484] = n_Body_y[484];
                c_Body_x[485] = n_Body_x[485];
                c_Body_y[485] = n_Body_y[485];
                c_Body_x[486] = n_Body_x[486];
                c_Body_y[486] = n_Body_y[486];
                c_Body_x[487] = n_Body_x[487];
                c_Body_y[487] = n_Body_y[487];
                c_Body_x[488] = n_Body_x[488];
                c_Body_y[488] = n_Body_y[488];
                c_Body_x[489] = n_Body_x[489];
                c_Body_y[489] = n_Body_y[489];
                c_Body_x[490] = n_Body_x[490];
                c_Body_y[490] = n_Body_y[490];
                c_Body_x[491] = n_Body_x[491];
                c_Body_y[491] = n_Body_y[491];
                c_Body_x[492] = n_Body_x[492];
                c_Body_y[492] = n_Body_y[492];
                c_Body_x[493] = n_Body_x[493];
                c_Body_y[493] = n_Body_y[493];
                c_Body_x[494] = n_Body_x[494];
                c_Body_y[494] = n_Body_y[494];
                c_Body_x[495] = n_Body_x[495];
                c_Body_y[495] = n_Body_y[495];
                c_Body_x[496] = n_Body_x[496];
                c_Body_y[496] = n_Body_y[496];
                c_Body_x[497] = n_Body_x[497];
                c_Body_y[497] = n_Body_y[497];
                c_Body_x[498] = n_Body_x[498];
                c_Body_y[498] = n_Body_y[498];
                c_Body_x[499] = n_Body_x[499];
                c_Body_y[499] = n_Body_y[499];
                c_Body_x[500] = n_Body_x[500];
                c_Body_y[500] = n_Body_y[500];
                c_Body_x[501] = n_Body_x[501];
                c_Body_y[501] = n_Body_y[501];
                c_Body_x[502] = n_Body_x[502];
                c_Body_y[502] = n_Body_y[502];
                c_Body_x[503] = n_Body_x[503];
                c_Body_y[503] = n_Body_y[503];
                c_Body_x[504] = n_Body_x[504];
                c_Body_y[504] = n_Body_y[504];
                c_Body_x[505] = n_Body_x[505];
                c_Body_y[505] = n_Body_y[505];
                c_Body_x[506] = n_Body_x[506];
                c_Body_y[506] = n_Body_y[506];
                c_Body_x[507] = n_Body_x[507];
                c_Body_y[507] = n_Body_y[507];
                c_Body_x[508] = n_Body_x[508];
                c_Body_y[508] = n_Body_y[508];
                c_Body_x[509] = n_Body_x[509];
                c_Body_y[509] = n_Body_y[509];
                c_Body_x[510] = n_Body_x[510];
                c_Body_y[510] = n_Body_y[510];
                c_Body_x[511] = n_Body_x[511];
                c_Body_y[511] = n_Body_y[511];
                c_Body_x[512] = n_Body_x[512];
                c_Body_y[512] = n_Body_y[512];
                c_Body_x[513] = n_Body_x[513];
                c_Body_y[513] = n_Body_y[513];
                c_Body_x[514] = n_Body_x[514];
                c_Body_y[514] = n_Body_y[514];
                c_Body_x[515] = n_Body_x[515];
                c_Body_y[515] = n_Body_y[515];
                c_Body_x[516] = n_Body_x[516];
                c_Body_y[516] = n_Body_y[516];
                c_Body_x[517] = n_Body_x[517];
                c_Body_y[517] = n_Body_y[517];
                c_Body_x[518] = n_Body_x[518];
                c_Body_y[518] = n_Body_y[518];
                c_Body_x[519] = n_Body_x[519];
                c_Body_y[519] = n_Body_y[519];
                c_Body_x[520] = n_Body_x[520];
                c_Body_y[520] = n_Body_y[520];
                c_Body_x[521] = n_Body_x[521];
                c_Body_y[521] = n_Body_y[521];
                c_Body_x[522] = n_Body_x[522];
                c_Body_y[522] = n_Body_y[522];
                c_Body_x[523] = n_Body_x[523];
                c_Body_y[523] = n_Body_y[523];
                c_Body_x[524] = n_Body_x[524];
                c_Body_y[524] = n_Body_y[524];
                c_Body_x[525] = n_Body_x[525];
                c_Body_y[525] = n_Body_y[525];
                c_Body_x[526] = n_Body_x[526];
                c_Body_y[526] = n_Body_y[526];
                c_Body_x[527] = n_Body_x[527];
                c_Body_y[527] = n_Body_y[527];
                c_Body_x[528] = n_Body_x[528];
                c_Body_y[528] = n_Body_y[528];
                c_Body_x[529] = n_Body_x[529];
                c_Body_y[529] = n_Body_y[529];
                c_Body_x[530] = n_Body_x[530];
                c_Body_y[530] = n_Body_y[530];
                c_Body_x[531] = n_Body_x[531];
                c_Body_y[531] = n_Body_y[531];
                c_Body_x[532] = n_Body_x[532];
                c_Body_y[532] = n_Body_y[532];
                c_Body_x[533] = n_Body_x[533];
                c_Body_y[533] = n_Body_y[533];
                c_Body_x[534] = n_Body_x[534];
                c_Body_y[534] = n_Body_y[534];
                c_Body_x[535] = n_Body_x[535];
                c_Body_y[535] = n_Body_y[535];
                c_Body_x[536] = n_Body_x[536];
                c_Body_y[536] = n_Body_y[536];
                c_Body_x[537] = n_Body_x[537];
                c_Body_y[537] = n_Body_y[537];
                c_Body_x[538] = n_Body_x[538];
                c_Body_y[538] = n_Body_y[538];
                c_Body_x[539] = n_Body_x[539];
                c_Body_y[539] = n_Body_y[539];
                c_Body_x[540] = n_Body_x[540];
                c_Body_y[540] = n_Body_y[540];
                c_Body_x[541] = n_Body_x[541];
                c_Body_y[541] = n_Body_y[541];
                c_Body_x[542] = n_Body_x[542];
                c_Body_y[542] = n_Body_y[542];
                c_Body_x[543] = n_Body_x[543];
                c_Body_y[543] = n_Body_y[543];
                c_Body_x[544] = n_Body_x[544];
                c_Body_y[544] = n_Body_y[544];
                c_Body_x[545] = n_Body_x[545];
                c_Body_y[545] = n_Body_y[545];
                c_Body_x[546] = n_Body_x[546];
                c_Body_y[546] = n_Body_y[546];
                c_Body_x[547] = n_Body_x[547];
                c_Body_y[547] = n_Body_y[547];
                c_Body_x[548] = n_Body_x[548];
                c_Body_y[548] = n_Body_y[548];
                c_Body_x[549] = n_Body_x[549];
                c_Body_y[549] = n_Body_y[549];
                c_Body_x[550] = n_Body_x[550];
                c_Body_y[550] = n_Body_y[550];
                c_Body_x[551] = n_Body_x[551];
                c_Body_y[551] = n_Body_y[551];
                c_Body_x[552] = n_Body_x[552];
                c_Body_y[552] = n_Body_y[552];
                c_Body_x[553] = n_Body_x[553];
                c_Body_y[553] = n_Body_y[553];
                c_Body_x[554] = n_Body_x[554];
                c_Body_y[554] = n_Body_y[554];
                c_Body_x[555] = n_Body_x[555];
                c_Body_y[555] = n_Body_y[555];
                c_Body_x[556] = n_Body_x[556];
                c_Body_y[556] = n_Body_y[556];
                c_Body_x[557] = n_Body_x[557];
                c_Body_y[557] = n_Body_y[557];
                c_Body_x[558] = n_Body_x[558];
                c_Body_y[558] = n_Body_y[558];
                c_Body_x[559] = n_Body_x[559];
                c_Body_y[559] = n_Body_y[559];
                c_Body_x[560] = n_Body_x[560];
                c_Body_y[560] = n_Body_y[560];
                c_Body_x[561] = n_Body_x[561];
                c_Body_y[561] = n_Body_y[561];
                c_Body_x[562] = n_Body_x[562];
                c_Body_y[562] = n_Body_y[562];
                c_Body_x[563] = n_Body_x[563];
                c_Body_y[563] = n_Body_y[563];
                c_Body_x[564] = n_Body_x[564];
                c_Body_y[564] = n_Body_y[564];
                c_Body_x[565] = n_Body_x[565];
                c_Body_y[565] = n_Body_y[565];
                c_Body_x[566] = n_Body_x[566];
                c_Body_y[566] = n_Body_y[566];
                c_Body_x[567] = n_Body_x[567];
                c_Body_y[567] = n_Body_y[567];
                c_Body_x[568] = n_Body_x[568];
                c_Body_y[568] = n_Body_y[568];
                c_Body_x[569] = n_Body_x[569];
                c_Body_y[569] = n_Body_y[569];
                c_Body_x[570] = n_Body_x[570];
                c_Body_y[570] = n_Body_y[570];
                c_Body_x[571] = n_Body_x[571];
                c_Body_y[571] = n_Body_y[571];
                c_Body_x[572] = n_Body_x[572];
                c_Body_y[572] = n_Body_y[572];
                c_Body_x[573] = n_Body_x[573];
                c_Body_y[573] = n_Body_y[573];
                c_Body_x[574] = n_Body_x[574];
                c_Body_y[574] = n_Body_y[574];
                c_Body_x[575] = n_Body_x[575];
                c_Body_y[575] = n_Body_y[575];
                c_Body_x[576] = n_Body_x[576];
                c_Body_y[576] = n_Body_y[576];
                c_Body_x[577] = n_Body_x[577];
                c_Body_y[577] = n_Body_y[577];
                c_Body_x[578] = n_Body_x[578];
                c_Body_y[578] = n_Body_y[578];
                c_Body_x[579] = n_Body_x[579];
                c_Body_y[579] = n_Body_y[579];
                c_Body_x[580] = n_Body_x[580];
                c_Body_y[580] = n_Body_y[580];
                c_Body_x[581] = n_Body_x[581];
                c_Body_y[581] = n_Body_y[581];
                c_Body_x[582] = n_Body_x[582];
                c_Body_y[582] = n_Body_y[582];
                c_Body_x[583] = n_Body_x[583];
                c_Body_y[583] = n_Body_y[583];
                c_Body_x[584] = n_Body_x[584];
                c_Body_y[584] = n_Body_y[584];
                c_Body_x[585] = n_Body_x[585];
                c_Body_y[585] = n_Body_y[585];
                c_Body_x[586] = n_Body_x[586];
                c_Body_y[586] = n_Body_y[586];
                c_Body_x[587] = n_Body_x[587];
                c_Body_y[587] = n_Body_y[587];
                c_Body_x[588] = n_Body_x[588];
                c_Body_y[588] = n_Body_y[588];
                c_Body_x[589] = n_Body_x[589];
                c_Body_y[589] = n_Body_y[589];
                c_Body_x[590] = n_Body_x[590];
                c_Body_y[590] = n_Body_y[590];
                c_Body_x[591] = n_Body_x[591];
                c_Body_y[591] = n_Body_y[591];
                c_Body_x[592] = n_Body_x[592];
                c_Body_y[592] = n_Body_y[592];
                c_Body_x[593] = n_Body_x[593];
                c_Body_y[593] = n_Body_y[593];
                c_Body_x[594] = n_Body_x[594];
                c_Body_y[594] = n_Body_y[594];
                c_Body_x[595] = n_Body_x[595];
                c_Body_y[595] = n_Body_y[595];
                c_Body_x[596] = n_Body_x[596];
                c_Body_y[596] = n_Body_y[596];
                c_Body_x[597] = n_Body_x[597];
                c_Body_y[597] = n_Body_y[597];
                c_Body_x[598] = n_Body_x[598];
                c_Body_y[598] = n_Body_y[598];
                c_Body_x[599] = n_Body_x[599];
                c_Body_y[599] = n_Body_y[599];
                c_Body_x[600] = n_Body_x[600];
                c_Body_y[600] = n_Body_y[600];
                c_Body_x[601] = n_Body_x[601];
                c_Body_y[601] = n_Body_y[601];
                c_Body_x[602] = n_Body_x[602];
                c_Body_y[602] = n_Body_y[602];
                c_Body_x[603] = n_Body_x[603];
                c_Body_y[603] = n_Body_y[603];
                c_Body_x[604] = n_Body_x[604];
                c_Body_y[604] = n_Body_y[604];
                c_Body_x[605] = n_Body_x[605];
                c_Body_y[605] = n_Body_y[605];
                c_Body_x[606] = n_Body_x[606];
                c_Body_y[606] = n_Body_y[606];
                c_Body_x[607] = n_Body_x[607];
                c_Body_y[607] = n_Body_y[607];
                c_Body_x[608] = n_Body_x[608];
                c_Body_y[608] = n_Body_y[608];
                c_Body_x[609] = n_Body_x[609];
                c_Body_y[609] = n_Body_y[609];
                c_Body_x[610] = n_Body_x[610];
                c_Body_y[610] = n_Body_y[610];
                c_Body_x[611] = n_Body_x[611];
                c_Body_y[611] = n_Body_y[611];
                c_Body_x[612] = n_Body_x[612];
                c_Body_y[612] = n_Body_y[612];
                c_Body_x[613] = n_Body_x[613];
                c_Body_y[613] = n_Body_y[613];
                c_Body_x[614] = n_Body_x[614];
                c_Body_y[614] = n_Body_y[614];
                c_Body_x[615] = n_Body_x[615];
                c_Body_y[615] = n_Body_y[615];
                c_Body_x[616] = n_Body_x[616];
                c_Body_y[616] = n_Body_y[616];
                c_Body_x[617] = n_Body_x[617];
                c_Body_y[617] = n_Body_y[617];
                c_Body_x[618] = n_Body_x[618];
                c_Body_y[618] = n_Body_y[618];
                c_Body_x[619] = n_Body_x[619];
                c_Body_y[619] = n_Body_y[619];
                c_Body_x[620] = n_Body_x[620];
                c_Body_y[620] = n_Body_y[620];
                c_Body_x[621] = n_Body_x[621];
                c_Body_y[621] = n_Body_y[621];
                c_Body_x[622] = n_Body_x[622];
                c_Body_y[622] = n_Body_y[622];
                c_Body_x[623] = n_Body_x[623];
                c_Body_y[623] = n_Body_y[623];
                c_Body_x[624] = n_Body_x[624];
                c_Body_y[624] = n_Body_y[624];
                c_Body_x[625] = n_Body_x[625];
                c_Body_y[625] = n_Body_y[625];
                c_Body_x[626] = n_Body_x[626];
                c_Body_y[626] = n_Body_y[626];
                c_Body_x[627] = n_Body_x[627];
                c_Body_y[627] = n_Body_y[627];
                c_Body_x[628] = n_Body_x[628];
                c_Body_y[628] = n_Body_y[628];
                c_Body_x[629] = n_Body_x[629];
                c_Body_y[629] = n_Body_y[629];
                c_Body_x[630] = n_Body_x[630];
                c_Body_y[630] = n_Body_y[630];
                c_Body_x[631] = n_Body_x[631];
                c_Body_y[631] = n_Body_y[631];
                c_Body_x[632] = n_Body_x[632];
                c_Body_y[632] = n_Body_y[632];
                c_Body_x[633] = n_Body_x[633];
                c_Body_y[633] = n_Body_y[633];
                c_Body_x[634] = n_Body_x[634];
                c_Body_y[634] = n_Body_y[634];
                c_Body_x[635] = n_Body_x[635];
                c_Body_y[635] = n_Body_y[635];
                c_Body_x[636] = n_Body_x[636];
                c_Body_y[636] = n_Body_y[636];
                c_Body_x[637] = n_Body_x[637];
                c_Body_y[637] = n_Body_y[637];
                c_Body_x[638] = n_Body_x[638];
                c_Body_y[638] = n_Body_y[638];
                c_Body_x[639] = n_Body_x[639];
                c_Body_y[639] = n_Body_y[639];
                c_Body_x[640] = n_Body_x[640];
                c_Body_y[640] = n_Body_y[640];
                c_Body_x[641] = n_Body_x[641];
                c_Body_y[641] = n_Body_y[641];
                c_Body_x[642] = n_Body_x[642];
                c_Body_y[642] = n_Body_y[642];
                c_Body_x[643] = n_Body_x[643];
                c_Body_y[643] = n_Body_y[643];
                c_Body_x[644] = n_Body_x[644];
                c_Body_y[644] = n_Body_y[644];
                c_Body_x[645] = n_Body_x[645];
                c_Body_y[645] = n_Body_y[645];
                c_Body_x[646] = n_Body_x[646];
                c_Body_y[646] = n_Body_y[646];
                c_Body_x[647] = n_Body_x[647];
                c_Body_y[647] = n_Body_y[647];
                c_Body_x[648] = n_Body_x[648];
                c_Body_y[648] = n_Body_y[648];
                c_Body_x[649] = n_Body_x[649];
                c_Body_y[649] = n_Body_y[649];
                c_Body_x[650] = n_Body_x[650];
                c_Body_y[650] = n_Body_y[650];
                c_Body_x[651] = n_Body_x[651];
                c_Body_y[651] = n_Body_y[651];
                c_Body_x[652] = n_Body_x[652];
                c_Body_y[652] = n_Body_y[652];
                c_Body_x[653] = n_Body_x[653];
                c_Body_y[653] = n_Body_y[653];
                c_Body_x[654] = n_Body_x[654];
                c_Body_y[654] = n_Body_y[654];
                c_Body_x[655] = n_Body_x[655];
                c_Body_y[655] = n_Body_y[655];
                c_Body_x[656] = n_Body_x[656];
                c_Body_y[656] = n_Body_y[656];
                c_Body_x[657] = n_Body_x[657];
                c_Body_y[657] = n_Body_y[657];
                c_Body_x[658] = n_Body_x[658];
                c_Body_y[658] = n_Body_y[658];
                c_Body_x[659] = n_Body_x[659];
                c_Body_y[659] = n_Body_y[659];
                c_Body_x[660] = n_Body_x[660];
                c_Body_y[660] = n_Body_y[660];
                c_Body_x[661] = n_Body_x[661];
                c_Body_y[661] = n_Body_y[661];
                c_Body_x[662] = n_Body_x[662];
                c_Body_y[662] = n_Body_y[662];
                c_Body_x[663] = n_Body_x[663];
                c_Body_y[663] = n_Body_y[663];
                c_Body_x[664] = n_Body_x[664];
                c_Body_y[664] = n_Body_y[664];
                c_Body_x[665] = n_Body_x[665];
                c_Body_y[665] = n_Body_y[665];
                c_Body_x[666] = n_Body_x[666];
                c_Body_y[666] = n_Body_y[666];
                c_Body_x[667] = n_Body_x[667];
                c_Body_y[667] = n_Body_y[667];
                c_Body_x[668] = n_Body_x[668];
                c_Body_y[668] = n_Body_y[668];
                c_Body_x[669] = n_Body_x[669];
                c_Body_y[669] = n_Body_y[669];
                c_Body_x[670] = n_Body_x[670];
                c_Body_y[670] = n_Body_y[670];
                c_Body_x[671] = n_Body_x[671];
                c_Body_y[671] = n_Body_y[671];
                c_Body_x[672] = n_Body_x[672];
                c_Body_y[672] = n_Body_y[672];
                c_Body_x[673] = n_Body_x[673];
                c_Body_y[673] = n_Body_y[673];
                c_Body_x[674] = n_Body_x[674];
                c_Body_y[674] = n_Body_y[674];
                c_Body_x[675] = n_Body_x[675];
                c_Body_y[675] = n_Body_y[675];
                c_Body_x[676] = n_Body_x[676];
                c_Body_y[676] = n_Body_y[676];
                c_Body_x[677] = n_Body_x[677];
                c_Body_y[677] = n_Body_y[677];
                c_Body_x[678] = n_Body_x[678];
                c_Body_y[678] = n_Body_y[678];
                c_Body_x[679] = n_Body_x[679];
                c_Body_y[679] = n_Body_y[679];
                c_Body_x[680] = n_Body_x[680];
                c_Body_y[680] = n_Body_y[680];
                c_Body_x[681] = n_Body_x[681];
                c_Body_y[681] = n_Body_y[681];
                c_Body_x[682] = n_Body_x[682];
                c_Body_y[682] = n_Body_y[682];
                c_Body_x[683] = n_Body_x[683];
                c_Body_y[683] = n_Body_y[683];
                c_Body_x[684] = n_Body_x[684];
                c_Body_y[684] = n_Body_y[684];
                c_Body_x[685] = n_Body_x[685];
                c_Body_y[685] = n_Body_y[685];
                c_Body_x[686] = n_Body_x[686];
                c_Body_y[686] = n_Body_y[686];
                c_Body_x[687] = n_Body_x[687];
                c_Body_y[687] = n_Body_y[687];
                c_Body_x[688] = n_Body_x[688];
                c_Body_y[688] = n_Body_y[688];
                c_Body_x[689] = n_Body_x[689];
                c_Body_y[689] = n_Body_y[689];
                c_Body_x[690] = n_Body_x[690];
                c_Body_y[690] = n_Body_y[690];
                c_Body_x[691] = n_Body_x[691];
                c_Body_y[691] = n_Body_y[691];
                c_Body_x[692] = n_Body_x[692];
                c_Body_y[692] = n_Body_y[692];
                c_Body_x[693] = n_Body_x[693];
                c_Body_y[693] = n_Body_y[693];
                c_Body_x[694] = n_Body_x[694];
                c_Body_y[694] = n_Body_y[694];
                c_Body_x[695] = n_Body_x[695];
                c_Body_y[695] = n_Body_y[695];
                c_Body_x[696] = n_Body_x[696];
                c_Body_y[696] = n_Body_y[696];
                c_Body_x[697] = n_Body_x[697];
                c_Body_y[697] = n_Body_y[697];
                c_Body_x[698] = n_Body_x[698];
                c_Body_y[698] = n_Body_y[698];
                c_Body_x[699] = n_Body_x[699];
                c_Body_y[699] = n_Body_y[699];
                c_Body_x[700] = n_Body_x[700];
                c_Body_y[700] = n_Body_y[700];
                c_Body_x[701] = n_Body_x[701];
                c_Body_y[701] = n_Body_y[701];
                c_Body_x[702] = n_Body_x[702];
                c_Body_y[702] = n_Body_y[702];
                c_Body_x[703] = n_Body_x[703];
                c_Body_y[703] = n_Body_y[703];
                c_Body_x[704] = n_Body_x[704];
                c_Body_y[704] = n_Body_y[704];
                c_Body_x[705] = n_Body_x[705];
                c_Body_y[705] = n_Body_y[705];
                c_Body_x[706] = n_Body_x[706];
                c_Body_y[706] = n_Body_y[706];
                c_Body_x[707] = n_Body_x[707];
                c_Body_y[707] = n_Body_y[707];
                c_Body_x[708] = n_Body_x[708];
                c_Body_y[708] = n_Body_y[708];
                c_Body_x[709] = n_Body_x[709];
                c_Body_y[709] = n_Body_y[709];
                c_Body_x[710] = n_Body_x[710];
                c_Body_y[710] = n_Body_y[710];
                c_Body_x[711] = n_Body_x[711];
                c_Body_y[711] = n_Body_y[711];
                c_Body_x[712] = n_Body_x[712];
                c_Body_y[712] = n_Body_y[712];
                c_Body_x[713] = n_Body_x[713];
                c_Body_y[713] = n_Body_y[713];
                c_Body_x[714] = n_Body_x[714];
                c_Body_y[714] = n_Body_y[714];
                c_Body_x[715] = n_Body_x[715];
                c_Body_y[715] = n_Body_y[715];
                c_Body_x[716] = n_Body_x[716];
                c_Body_y[716] = n_Body_y[716];
                c_Body_x[717] = n_Body_x[717];
                c_Body_y[717] = n_Body_y[717];
                c_Body_x[718] = n_Body_x[718];
                c_Body_y[718] = n_Body_y[718];
                c_Body_x[719] = n_Body_x[719];
                c_Body_y[719] = n_Body_y[719];
                c_Body_x[720] = n_Body_x[720];
                c_Body_y[720] = n_Body_y[720];
                c_Body_x[721] = n_Body_x[721];
                c_Body_y[721] = n_Body_y[721];
                c_Body_x[722] = n_Body_x[722];
                c_Body_y[722] = n_Body_y[722];
                c_Body_x[723] = n_Body_x[723];
                c_Body_y[723] = n_Body_y[723];
                c_Body_x[724] = n_Body_x[724];
                c_Body_y[724] = n_Body_y[724];
                c_Body_x[725] = n_Body_x[725];
                c_Body_y[725] = n_Body_y[725];
                c_Body_x[726] = n_Body_x[726];
                c_Body_y[726] = n_Body_y[726];
                c_Body_x[727] = n_Body_x[727];
                c_Body_y[727] = n_Body_y[727];
                c_Body_x[728] = n_Body_x[728];
                c_Body_y[728] = n_Body_y[728];
                c_Body_x[729] = n_Body_x[729];
                c_Body_y[729] = n_Body_y[729];
                c_Body_x[730] = n_Body_x[730];
                c_Body_y[730] = n_Body_y[730];
                c_Body_x[731] = n_Body_x[731];
                c_Body_y[731] = n_Body_y[731];
                c_Body_x[732] = n_Body_x[732];
                c_Body_y[732] = n_Body_y[732];
                c_Body_x[733] = n_Body_x[733];
                c_Body_y[733] = n_Body_y[733];
                c_Body_x[734] = n_Body_x[734];
                c_Body_y[734] = n_Body_y[734];
                c_Body_x[735] = n_Body_x[735];
                c_Body_y[735] = n_Body_y[735];
                c_Body_x[736] = n_Body_x[736];
                c_Body_y[736] = n_Body_y[736];
                c_Body_x[737] = n_Body_x[737];
                c_Body_y[737] = n_Body_y[737];
                c_Body_x[738] = n_Body_x[738];
                c_Body_y[738] = n_Body_y[738];
                c_Body_x[739] = n_Body_x[739];
                c_Body_y[739] = n_Body_y[739];
                c_Body_x[740] = n_Body_x[740];
                c_Body_y[740] = n_Body_y[740];
                c_Body_x[741] = n_Body_x[741];
                c_Body_y[741] = n_Body_y[741];
                c_Body_x[742] = n_Body_x[742];
                c_Body_y[742] = n_Body_y[742];
                c_Body_x[743] = n_Body_x[743];
                c_Body_y[743] = n_Body_y[743];
                c_Body_x[744] = n_Body_x[744];
                c_Body_y[744] = n_Body_y[744];
                c_Body_x[745] = n_Body_x[745];
                c_Body_y[745] = n_Body_y[745];
                c_Body_x[746] = n_Body_x[746];
                c_Body_y[746] = n_Body_y[746];
                c_Body_x[747] = n_Body_x[747];
                c_Body_y[747] = n_Body_y[747];
                c_Body_x[748] = n_Body_x[748];
                c_Body_y[748] = n_Body_y[748];
                c_Body_x[749] = n_Body_x[749];
                c_Body_y[749] = n_Body_y[749];
                c_Body_x[750] = n_Body_x[750];
                c_Body_y[750] = n_Body_y[750];
                c_Body_x[751] = n_Body_x[751];
                c_Body_y[751] = n_Body_y[751];
                c_Body_x[752] = n_Body_x[752];
                c_Body_y[752] = n_Body_y[752];
                c_Body_x[753] = n_Body_x[753];
                c_Body_y[753] = n_Body_y[753];
                c_Body_x[754] = n_Body_x[754];
                c_Body_y[754] = n_Body_y[754];
                c_Body_x[755] = n_Body_x[755];
                c_Body_y[755] = n_Body_y[755];
                c_Body_x[756] = n_Body_x[756];
                c_Body_y[756] = n_Body_y[756];
                c_Body_x[757] = n_Body_x[757];
                c_Body_y[757] = n_Body_y[757];
                c_Body_x[758] = n_Body_x[758];
                c_Body_y[758] = n_Body_y[758];
                c_Body_x[759] = n_Body_x[759];
                c_Body_y[759] = n_Body_y[759];
                c_Body_x[760] = n_Body_x[760];
                c_Body_y[760] = n_Body_y[760];
                c_Body_x[761] = n_Body_x[761];
                c_Body_y[761] = n_Body_y[761];
                c_Body_x[762] = n_Body_x[762];
                c_Body_y[762] = n_Body_y[762];
                c_Body_x[763] = n_Body_x[763];
                c_Body_y[763] = n_Body_y[763];
                c_Body_x[764] = n_Body_x[764];
                c_Body_y[764] = n_Body_y[764];
                c_Body_x[765] = n_Body_x[765];
                c_Body_y[765] = n_Body_y[765];
                c_Body_x[766] = n_Body_x[766];
                c_Body_y[766] = n_Body_y[766];
                c_Body_x[767] = n_Body_x[767];
                c_Body_y[767] = n_Body_y[767];
                c_Body_x[768] = n_Body_x[768];
                c_Body_y[768] = n_Body_y[768];
                c_Body_x[769] = n_Body_x[769];
                c_Body_y[769] = n_Body_y[769];
                c_Body_x[770] = n_Body_x[770];
                c_Body_y[770] = n_Body_y[770];
                c_Body_x[771] = n_Body_x[771];
                c_Body_y[771] = n_Body_y[771];
                c_Body_x[772] = n_Body_x[772];
                c_Body_y[772] = n_Body_y[772];
                c_Body_x[773] = n_Body_x[773];
                c_Body_y[773] = n_Body_y[773];
                c_Body_x[774] = n_Body_x[774];
                c_Body_y[774] = n_Body_y[774];
                c_Body_x[775] = n_Body_x[775];
                c_Body_y[775] = n_Body_y[775];
                c_Body_x[776] = n_Body_x[776];
                c_Body_y[776] = n_Body_y[776];
                c_Body_x[777] = n_Body_x[777];
                c_Body_y[777] = n_Body_y[777];
                c_Body_x[778] = n_Body_x[778];
                c_Body_y[778] = n_Body_y[778];
                c_Body_x[779] = n_Body_x[779];
                c_Body_y[779] = n_Body_y[779];
                c_Body_x[780] = n_Body_x[780];
                c_Body_y[780] = n_Body_y[780];
                c_Body_x[781] = n_Body_x[781];
                c_Body_y[781] = n_Body_y[781];
                c_Body_x[782] = n_Body_x[782];
                c_Body_y[782] = n_Body_y[782];
                c_Body_x[783] = n_Body_x[783];
                c_Body_y[783] = n_Body_y[783];
                c_Body_x[784] = n_Body_x[784];
                c_Body_y[784] = n_Body_y[784];
                c_Body_x[785] = n_Body_x[785];
                c_Body_y[785] = n_Body_y[785];
                c_Body_x[786] = n_Body_x[786];
                c_Body_y[786] = n_Body_y[786];
                c_Body_x[787] = n_Body_x[787];
                c_Body_y[787] = n_Body_y[787];
                c_Body_x[788] = n_Body_x[788];
                c_Body_y[788] = n_Body_y[788];
                c_Body_x[789] = n_Body_x[789];
                c_Body_y[789] = n_Body_y[789];
                c_Body_x[790] = n_Body_x[790];
                c_Body_y[790] = n_Body_y[790];
                c_Body_x[791] = n_Body_x[791];
                c_Body_y[791] = n_Body_y[791];
                c_Body_x[792] = n_Body_x[792];
                c_Body_y[792] = n_Body_y[792];
                c_Body_x[793] = n_Body_x[793];
                c_Body_y[793] = n_Body_y[793];
                c_Body_x[794] = n_Body_x[794];
                c_Body_y[794] = n_Body_y[794];
                c_Body_x[795] = n_Body_x[795];
                c_Body_y[795] = n_Body_y[795];
                c_Body_x[796] = n_Body_x[796];
                c_Body_y[796] = n_Body_y[796];
                c_Body_x[797] = n_Body_x[797];
                c_Body_y[797] = n_Body_y[797];
                c_Body_x[798] = n_Body_x[798];
                c_Body_y[798] = n_Body_y[798];
                c_Body_x[799] = n_Body_x[799];
                c_Body_y[799] = n_Body_y[799];
                c_Body_x[800] = n_Body_x[800];
                c_Body_y[800] = n_Body_y[800];
                c_Body_x[801] = n_Body_x[801];
                c_Body_y[801] = n_Body_y[801];
                c_Body_x[802] = n_Body_x[802];
                c_Body_y[802] = n_Body_y[802];
                c_Body_x[803] = n_Body_x[803];
                c_Body_y[803] = n_Body_y[803];
                c_Body_x[804] = n_Body_x[804];
                c_Body_y[804] = n_Body_y[804];
                c_Body_x[805] = n_Body_x[805];
                c_Body_y[805] = n_Body_y[805];
                c_Body_x[806] = n_Body_x[806];
                c_Body_y[806] = n_Body_y[806];
                c_Body_x[807] = n_Body_x[807];
                c_Body_y[807] = n_Body_y[807];
                c_Body_x[808] = n_Body_x[808];
                c_Body_y[808] = n_Body_y[808];
                c_Body_x[809] = n_Body_x[809];
                c_Body_y[809] = n_Body_y[809];
                c_Body_x[810] = n_Body_x[810];
                c_Body_y[810] = n_Body_y[810];
                c_Body_x[811] = n_Body_x[811];
                c_Body_y[811] = n_Body_y[811];
                c_Body_x[812] = n_Body_x[812];
                c_Body_y[812] = n_Body_y[812];
                c_Body_x[813] = n_Body_x[813];
                c_Body_y[813] = n_Body_y[813];
                c_Body_x[814] = n_Body_x[814];
                c_Body_y[814] = n_Body_y[814];
                c_Body_x[815] = n_Body_x[815];
                c_Body_y[815] = n_Body_y[815];
                c_Body_x[816] = n_Body_x[816];
                c_Body_y[816] = n_Body_y[816];
                c_Body_x[817] = n_Body_x[817];
                c_Body_y[817] = n_Body_y[817];
                c_Body_x[818] = n_Body_x[818];
                c_Body_y[818] = n_Body_y[818];
                c_Body_x[819] = n_Body_x[819];
                c_Body_y[819] = n_Body_y[819];
                c_Body_x[820] = n_Body_x[820];
                c_Body_y[820] = n_Body_y[820];
                c_Body_x[821] = n_Body_x[821];
                c_Body_y[821] = n_Body_y[821];
                c_Body_x[822] = n_Body_x[822];
                c_Body_y[822] = n_Body_y[822];
                c_Body_x[823] = n_Body_x[823];
                c_Body_y[823] = n_Body_y[823];
                c_Body_x[824] = n_Body_x[824];
                c_Body_y[824] = n_Body_y[824];
                c_Body_x[825] = n_Body_x[825];
                c_Body_y[825] = n_Body_y[825];
                c_Body_x[826] = n_Body_x[826];
                c_Body_y[826] = n_Body_y[826];
                c_Body_x[827] = n_Body_x[827];
                c_Body_y[827] = n_Body_y[827];
                c_Body_x[828] = n_Body_x[828];
                c_Body_y[828] = n_Body_y[828];
                c_Body_x[829] = n_Body_x[829];
                c_Body_y[829] = n_Body_y[829];
                c_Body_x[830] = n_Body_x[830];
                c_Body_y[830] = n_Body_y[830];
                c_Body_x[831] = n_Body_x[831];
                c_Body_y[831] = n_Body_y[831];
                c_Body_x[832] = n_Body_x[832];
                c_Body_y[832] = n_Body_y[832];
                c_Body_x[833] = n_Body_x[833];
                c_Body_y[833] = n_Body_y[833];
                c_Body_x[834] = n_Body_x[834];
                c_Body_y[834] = n_Body_y[834];
                c_Body_x[835] = n_Body_x[835];
                c_Body_y[835] = n_Body_y[835];
                c_Body_x[836] = n_Body_x[836];
                c_Body_y[836] = n_Body_y[836];
                c_Body_x[837] = n_Body_x[837];
                c_Body_y[837] = n_Body_y[837];
                c_Body_x[838] = n_Body_x[838];
                c_Body_y[838] = n_Body_y[838];
                c_Body_x[839] = n_Body_x[839];
                c_Body_y[839] = n_Body_y[839];
                c_Body_x[840] = n_Body_x[840];
                c_Body_y[840] = n_Body_y[840];
                c_Body_x[841] = n_Body_x[841];
                c_Body_y[841] = n_Body_y[841];
                c_Body_x[842] = n_Body_x[842];
                c_Body_y[842] = n_Body_y[842];
                c_Body_x[843] = n_Body_x[843];
                c_Body_y[843] = n_Body_y[843];
                c_Body_x[844] = n_Body_x[844];
                c_Body_y[844] = n_Body_y[844];
                c_Body_x[845] = n_Body_x[845];
                c_Body_y[845] = n_Body_y[845];
                c_Body_x[846] = n_Body_x[846];
                c_Body_y[846] = n_Body_y[846];
                c_Body_x[847] = n_Body_x[847];
                c_Body_y[847] = n_Body_y[847];
                c_Body_x[848] = n_Body_x[848];
                c_Body_y[848] = n_Body_y[848];
                c_Body_x[849] = n_Body_x[849];
                c_Body_y[849] = n_Body_y[849];
                c_Body_x[850] = n_Body_x[850];
                c_Body_y[850] = n_Body_y[850];
                c_Body_x[851] = n_Body_x[851];
                c_Body_y[851] = n_Body_y[851];
                c_Body_x[852] = n_Body_x[852];
                c_Body_y[852] = n_Body_y[852];
                c_Body_x[853] = n_Body_x[853];
                c_Body_y[853] = n_Body_y[853];
                c_Body_x[854] = n_Body_x[854];
                c_Body_y[854] = n_Body_y[854];
                c_Body_x[855] = n_Body_x[855];
                c_Body_y[855] = n_Body_y[855];
                c_Body_x[856] = n_Body_x[856];
                c_Body_y[856] = n_Body_y[856];
                c_Body_x[857] = n_Body_x[857];
                c_Body_y[857] = n_Body_y[857];
                c_Body_x[858] = n_Body_x[858];
                c_Body_y[858] = n_Body_y[858];
                c_Body_x[859] = n_Body_x[859];
                c_Body_y[859] = n_Body_y[859];
                c_Body_x[860] = n_Body_x[860];
                c_Body_y[860] = n_Body_y[860];
                c_Body_x[861] = n_Body_x[861];
                c_Body_y[861] = n_Body_y[861];
                c_Body_x[862] = n_Body_x[862];
                c_Body_y[862] = n_Body_y[862];
                c_Body_x[863] = n_Body_x[863];
                c_Body_y[863] = n_Body_y[863];
                c_Body_x[864] = n_Body_x[864];
                c_Body_y[864] = n_Body_y[864];
                c_Body_x[865] = n_Body_x[865];
                c_Body_y[865] = n_Body_y[865];
                c_Body_x[866] = n_Body_x[866];
                c_Body_y[866] = n_Body_y[866];
                c_Body_x[867] = n_Body_x[867];
                c_Body_y[867] = n_Body_y[867];
                c_Body_x[868] = n_Body_x[868];
                c_Body_y[868] = n_Body_y[868];
                c_Body_x[869] = n_Body_x[869];
                c_Body_y[869] = n_Body_y[869];
                c_Body_x[870] = n_Body_x[870];
                c_Body_y[870] = n_Body_y[870];
                c_Body_x[871] = n_Body_x[871];
                c_Body_y[871] = n_Body_y[871];
                c_Body_x[872] = n_Body_x[872];
                c_Body_y[872] = n_Body_y[872];
                c_Body_x[873] = n_Body_x[873];
                c_Body_y[873] = n_Body_y[873];
                c_Body_x[874] = n_Body_x[874];
                c_Body_y[874] = n_Body_y[874];
                c_Body_x[875] = n_Body_x[875];
                c_Body_y[875] = n_Body_y[875];
                c_Body_x[876] = n_Body_x[876];
                c_Body_y[876] = n_Body_y[876];
                c_Body_x[877] = n_Body_x[877];
                c_Body_y[877] = n_Body_y[877];
                c_Body_x[878] = n_Body_x[878];
                c_Body_y[878] = n_Body_y[878];
                c_Body_x[879] = n_Body_x[879];
                c_Body_y[879] = n_Body_y[879];
                c_Body_x[880] = n_Body_x[880];
                c_Body_y[880] = n_Body_y[880];
                c_Body_x[881] = n_Body_x[881];
                c_Body_y[881] = n_Body_y[881];
                c_Body_x[882] = n_Body_x[882];
                c_Body_y[882] = n_Body_y[882];
                c_Body_x[883] = n_Body_x[883];
                c_Body_y[883] = n_Body_y[883];
                c_Body_x[884] = n_Body_x[884];
                c_Body_y[884] = n_Body_y[884];
                c_Body_x[885] = n_Body_x[885];
                c_Body_y[885] = n_Body_y[885];
                c_Body_x[886] = n_Body_x[886];
                c_Body_y[886] = n_Body_y[886];
                c_Body_x[887] = n_Body_x[887];
                c_Body_y[887] = n_Body_y[887];
                c_Body_x[888] = n_Body_x[888];
                c_Body_y[888] = n_Body_y[888];
                c_Body_x[889] = n_Body_x[889];
                c_Body_y[889] = n_Body_y[889];
                c_Body_x[890] = n_Body_x[890];
                c_Body_y[890] = n_Body_y[890];
                c_Body_x[891] = n_Body_x[891];
                c_Body_y[891] = n_Body_y[891];
                c_Body_x[892] = n_Body_x[892];
                c_Body_y[892] = n_Body_y[892];
                c_Body_x[893] = n_Body_x[893];
                c_Body_y[893] = n_Body_y[893];
                c_Body_x[894] = n_Body_x[894];
                c_Body_y[894] = n_Body_y[894];
                c_Body_x[895] = n_Body_x[895];
                c_Body_y[895] = n_Body_y[895];
                c_Body_x[896] = n_Body_x[896];
                c_Body_y[896] = n_Body_y[896];
                c_Body_x[897] = n_Body_x[897];
                c_Body_y[897] = n_Body_y[897];
                c_Body_x[898] = n_Body_x[898];
                c_Body_y[898] = n_Body_y[898];
                c_Body_x[899] = n_Body_x[899];
                c_Body_y[899] = n_Body_y[899];
                c_Body_x[900] = n_Body_x[900];
                c_Body_y[900] = n_Body_y[900];
                c_Body_x[901] = n_Body_x[901];
                c_Body_y[901] = n_Body_y[901];
                c_Body_x[902] = n_Body_x[902];
                c_Body_y[902] = n_Body_y[902];
                c_Body_x[903] = n_Body_x[903];
                c_Body_y[903] = n_Body_y[903];
                c_Body_x[904] = n_Body_x[904];
                c_Body_y[904] = n_Body_y[904];
                c_Body_x[905] = n_Body_x[905];
                c_Body_y[905] = n_Body_y[905];
                c_Body_x[906] = n_Body_x[906];
                c_Body_y[906] = n_Body_y[906];
                c_Body_x[907] = n_Body_x[907];
                c_Body_y[907] = n_Body_y[907];
                c_Body_x[908] = n_Body_x[908];
                c_Body_y[908] = n_Body_y[908];
                c_Body_x[909] = n_Body_x[909];
                c_Body_y[909] = n_Body_y[909];
                c_Body_x[910] = n_Body_x[910];
                c_Body_y[910] = n_Body_y[910];
                c_Body_x[911] = n_Body_x[911];
                c_Body_y[911] = n_Body_y[911];
                c_Body_x[912] = n_Body_x[912];
                c_Body_y[912] = n_Body_y[912];
                c_Body_x[913] = n_Body_x[913];
                c_Body_y[913] = n_Body_y[913];
                c_Body_x[914] = n_Body_x[914];
                c_Body_y[914] = n_Body_y[914];
                c_Body_x[915] = n_Body_x[915];
                c_Body_y[915] = n_Body_y[915];
                c_Body_x[916] = n_Body_x[916];
                c_Body_y[916] = n_Body_y[916];
                c_Body_x[917] = n_Body_x[917];
                c_Body_y[917] = n_Body_y[917];
                c_Body_x[918] = n_Body_x[918];
                c_Body_y[918] = n_Body_y[918];
                c_Body_x[919] = n_Body_x[919];
                c_Body_y[919] = n_Body_y[919];
                c_Body_x[920] = n_Body_x[920];
                c_Body_y[920] = n_Body_y[920];
                c_Body_x[921] = n_Body_x[921];
                c_Body_y[921] = n_Body_y[921];
                c_Body_x[922] = n_Body_x[922];
                c_Body_y[922] = n_Body_y[922];
                c_Body_x[923] = n_Body_x[923];
                c_Body_y[923] = n_Body_y[923];
                c_Body_x[924] = n_Body_x[924];
                c_Body_y[924] = n_Body_y[924];
                c_Body_x[925] = n_Body_x[925];
                c_Body_y[925] = n_Body_y[925];
                c_Body_x[926] = n_Body_x[926];
                c_Body_y[926] = n_Body_y[926];
                c_Body_x[927] = n_Body_x[927];
                c_Body_y[927] = n_Body_y[927];
                c_Body_x[928] = n_Body_x[928];
                c_Body_y[928] = n_Body_y[928];
                c_Body_x[929] = n_Body_x[929];
                c_Body_y[929] = n_Body_y[929];
                c_Body_x[930] = n_Body_x[930];
                c_Body_y[930] = n_Body_y[930];
                c_Body_x[931] = n_Body_x[931];
                c_Body_y[931] = n_Body_y[931];
                c_Body_x[932] = n_Body_x[932];
                c_Body_y[932] = n_Body_y[932];
                c_Body_x[933] = n_Body_x[933];
                c_Body_y[933] = n_Body_y[933];
                c_Body_x[934] = n_Body_x[934];
                c_Body_y[934] = n_Body_y[934];
                c_Body_x[935] = n_Body_x[935];
                c_Body_y[935] = n_Body_y[935];
                c_Body_x[936] = n_Body_x[936];
                c_Body_y[936] = n_Body_y[936];
                c_Body_x[937] = n_Body_x[937];
                c_Body_y[937] = n_Body_y[937];
                c_Body_x[938] = n_Body_x[938];
                c_Body_y[938] = n_Body_y[938];
                c_Body_x[939] = n_Body_x[939];
                c_Body_y[939] = n_Body_y[939];
                c_Body_x[940] = n_Body_x[940];
                c_Body_y[940] = n_Body_y[940];
                c_Body_x[941] = n_Body_x[941];
                c_Body_y[941] = n_Body_y[941];
                c_Body_x[942] = n_Body_x[942];
                c_Body_y[942] = n_Body_y[942];
                c_Body_x[943] = n_Body_x[943];
                c_Body_y[943] = n_Body_y[943];
                c_Body_x[944] = n_Body_x[944];
                c_Body_y[944] = n_Body_y[944];
                c_Body_x[945] = n_Body_x[945];
                c_Body_y[945] = n_Body_y[945];
                c_Body_x[946] = n_Body_x[946];
                c_Body_y[946] = n_Body_y[946];
                c_Body_x[947] = n_Body_x[947];
                c_Body_y[947] = n_Body_y[947];
                c_Body_x[948] = n_Body_x[948];
                c_Body_y[948] = n_Body_y[948];
                c_Body_x[949] = n_Body_x[949];
                c_Body_y[949] = n_Body_y[949];
                c_Body_x[950] = n_Body_x[950];
                c_Body_y[950] = n_Body_y[950];
                c_Body_x[951] = n_Body_x[951];
                c_Body_y[951] = n_Body_y[951];
                c_Body_x[952] = n_Body_x[952];
                c_Body_y[952] = n_Body_y[952];
                c_Body_x[953] = n_Body_x[953];
                c_Body_y[953] = n_Body_y[953];
                c_Body_x[954] = n_Body_x[954];
                c_Body_y[954] = n_Body_y[954];
                c_Body_x[955] = n_Body_x[955];
                c_Body_y[955] = n_Body_y[955];
                c_Body_x[956] = n_Body_x[956];
                c_Body_y[956] = n_Body_y[956];
                c_Body_x[957] = n_Body_x[957];
                c_Body_y[957] = n_Body_y[957];
                c_Body_x[958] = n_Body_x[958];
                c_Body_y[958] = n_Body_y[958];
                c_Body_x[959] = n_Body_x[959];
                c_Body_y[959] = n_Body_y[959];
                c_Body_x[960] = n_Body_x[960];
                c_Body_y[960] = n_Body_y[960];
                c_Body_x[961] = n_Body_x[961];
                c_Body_y[961] = n_Body_y[961];
                c_Body_x[962] = n_Body_x[962];
                c_Body_y[962] = n_Body_y[962];
                c_Body_x[963] = n_Body_x[963];
                c_Body_y[963] = n_Body_y[963];
                c_Body_x[964] = n_Body_x[964];
                c_Body_y[964] = n_Body_y[964];
                c_Body_x[965] = n_Body_x[965];
                c_Body_y[965] = n_Body_y[965];
                c_Body_x[966] = n_Body_x[966];
                c_Body_y[966] = n_Body_y[966];
                c_Body_x[967] = n_Body_x[967];
                c_Body_y[967] = n_Body_y[967];
                c_Body_x[968] = n_Body_x[968];
                c_Body_y[968] = n_Body_y[968];
                c_Body_x[969] = n_Body_x[969];
                c_Body_y[969] = n_Body_y[969];
                c_Body_x[970] = n_Body_x[970];
                c_Body_y[970] = n_Body_y[970];
                c_Body_x[971] = n_Body_x[971];
                c_Body_y[971] = n_Body_y[971];
                c_Body_x[972] = n_Body_x[972];
                c_Body_y[972] = n_Body_y[972];
                c_Body_x[973] = n_Body_x[973];
                c_Body_y[973] = n_Body_y[973];
                c_Body_x[974] = n_Body_x[974];
                c_Body_y[974] = n_Body_y[974];
                c_Body_x[975] = n_Body_x[975];
                c_Body_y[975] = n_Body_y[975];
                c_Body_x[976] = n_Body_x[976];
                c_Body_y[976] = n_Body_y[976];
                c_Body_x[977] = n_Body_x[977];
                c_Body_y[977] = n_Body_y[977];
                c_Body_x[978] = n_Body_x[978];
                c_Body_y[978] = n_Body_y[978];
                c_Body_x[979] = n_Body_x[979];
                c_Body_y[979] = n_Body_y[979];
                c_Body_x[980] = n_Body_x[980];
                c_Body_y[980] = n_Body_y[980];
                c_Body_x[981] = n_Body_x[981];
                c_Body_y[981] = n_Body_y[981];
                c_Body_x[982] = n_Body_x[982];
                c_Body_y[982] = n_Body_y[982];
                c_Body_x[983] = n_Body_x[983];
                c_Body_y[983] = n_Body_y[983];
                c_Body_x[984] = n_Body_x[984];
                c_Body_y[984] = n_Body_y[984];
                c_Body_x[985] = n_Body_x[985];
                c_Body_y[985] = n_Body_y[985];
                c_Body_x[986] = n_Body_x[986];
                c_Body_y[986] = n_Body_y[986];
                c_Body_x[987] = n_Body_x[987];
                c_Body_y[987] = n_Body_y[987];
                c_Body_x[988] = n_Body_x[988];
                c_Body_y[988] = n_Body_y[988];
                c_Body_x[989] = n_Body_x[989];
                c_Body_y[989] = n_Body_y[989];
                c_Body_x[990] = n_Body_x[990];
                c_Body_y[990] = n_Body_y[990];
                c_Body_x[991] = n_Body_x[991];
                c_Body_y[991] = n_Body_y[991];
                c_Body_x[992] = n_Body_x[992];
                c_Body_y[992] = n_Body_y[992];
                c_Body_x[993] = n_Body_x[993];
                c_Body_y[993] = n_Body_y[993];
                c_Body_x[994] = n_Body_x[994];
                c_Body_y[994] = n_Body_y[994];
                c_Body_x[995] = n_Body_x[995];
                c_Body_y[995] = n_Body_y[995];
                c_Body_x[996] = n_Body_x[996];
                c_Body_y[996] = n_Body_y[996];
                c_Body_x[997] = n_Body_x[997];
                c_Body_y[997] = n_Body_y[997];
                c_Body_x[998] = n_Body_x[998];
                c_Body_y[998] = n_Body_y[998];
                c_Body_x[999] = n_Body_x[999];
                c_Body_y[999] = n_Body_y[999];
                c_Body_x[1000] = n_Body_x[1000];
                c_Body_y[1000] = n_Body_y[1000];
                c_Body_x[1001] = n_Body_x[1001];
                c_Body_y[1001] = n_Body_y[1001];
                c_Body_x[1002] = n_Body_x[1002];
                c_Body_y[1002] = n_Body_y[1002];
                c_Body_x[1003] = n_Body_x[1003];
                c_Body_y[1003] = n_Body_y[1003];
                c_Body_x[1004] = n_Body_x[1004];
                c_Body_y[1004] = n_Body_y[1004];
                c_Body_x[1005] = n_Body_x[1005];
                c_Body_y[1005] = n_Body_y[1005];
                c_Body_x[1006] = n_Body_x[1006];
                c_Body_y[1006] = n_Body_y[1006];
                c_Body_x[1007] = n_Body_x[1007];
                c_Body_y[1007] = n_Body_y[1007];
                c_Body_x[1008] = n_Body_x[1008];
                c_Body_y[1008] = n_Body_y[1008];
                c_Body_x[1009] = n_Body_x[1009];
                c_Body_y[1009] = n_Body_y[1009];
                c_Body_x[1010] = n_Body_x[1010];
                c_Body_y[1010] = n_Body_y[1010];
                c_Body_x[1011] = n_Body_x[1011];
                c_Body_y[1011] = n_Body_y[1011];
                c_Body_x[1012] = n_Body_x[1012];
                c_Body_y[1012] = n_Body_y[1012];
                c_Body_x[1013] = n_Body_x[1013];
                c_Body_y[1013] = n_Body_y[1013];
                c_Body_x[1014] = n_Body_x[1014];
                c_Body_y[1014] = n_Body_y[1014];
                c_Body_x[1015] = n_Body_x[1015];
                c_Body_y[1015] = n_Body_y[1015];
                c_Body_x[1016] = n_Body_x[1016];
                c_Body_y[1016] = n_Body_y[1016];
                c_Body_x[1017] = n_Body_x[1017];
                c_Body_y[1017] = n_Body_y[1017];
                c_Body_x[1018] = n_Body_x[1018];
                c_Body_y[1018] = n_Body_y[1018];
                c_Body_x[1019] = n_Body_x[1019];
                c_Body_y[1019] = n_Body_y[1019];
                c_Body_x[1020] = n_Body_x[1020];
                c_Body_y[1020] = n_Body_y[1020];
                c_Body_x[1021] = n_Body_x[1021];
                c_Body_y[1021] = n_Body_y[1021];
                c_Body_x[1022] = n_Body_x[1022];
                c_Body_y[1022] = n_Body_y[1022];
                c_Body_x[1023] = n_Body_x[1023];
                c_Body_y[1023] = n_Body_y[1023];
                c_Body_x[1024] = n_Body_x[1024];
                c_Body_y[1024] = n_Body_y[1024];
                c_Body_x[1025] = n_Body_x[1025];
                c_Body_y[1025] = n_Body_y[1025];
                c_Body_x[1026] = n_Body_x[1026];
                c_Body_y[1026] = n_Body_y[1026];
                c_Body_x[1027] = n_Body_x[1027];
                c_Body_y[1027] = n_Body_y[1027];
                c_Body_x[1028] = n_Body_x[1028];
                c_Body_y[1028] = n_Body_y[1028];
                c_Body_x[1029] = n_Body_x[1029];
                c_Body_y[1029] = n_Body_y[1029];
                c_Body_x[1030] = n_Body_x[1030];
                c_Body_y[1030] = n_Body_y[1030];
                c_Body_x[1031] = n_Body_x[1031];
                c_Body_y[1031] = n_Body_y[1031];
                c_Body_x[1032] = n_Body_x[1032];
                c_Body_y[1032] = n_Body_y[1032];
                c_Body_x[1033] = n_Body_x[1033];
                c_Body_y[1033] = n_Body_y[1033];
                c_Body_x[1034] = n_Body_x[1034];
                c_Body_y[1034] = n_Body_y[1034];
                c_Body_x[1035] = n_Body_x[1035];
                c_Body_y[1035] = n_Body_y[1035];
                c_Body_x[1036] = n_Body_x[1036];
                c_Body_y[1036] = n_Body_y[1036];
                c_Body_x[1037] = n_Body_x[1037];
                c_Body_y[1037] = n_Body_y[1037];
                c_Body_x[1038] = n_Body_x[1038];
                c_Body_y[1038] = n_Body_y[1038];
                c_Body_x[1039] = n_Body_x[1039];
                c_Body_y[1039] = n_Body_y[1039];
                c_Body_x[1040] = n_Body_x[1040];
                c_Body_y[1040] = n_Body_y[1040];
                c_Body_x[1041] = n_Body_x[1041];
                c_Body_y[1041] = n_Body_y[1041];
                c_Body_x[1042] = n_Body_x[1042];
                c_Body_y[1042] = n_Body_y[1042];
                c_Body_x[1043] = n_Body_x[1043];
                c_Body_y[1043] = n_Body_y[1043];
                c_Body_x[1044] = n_Body_x[1044];
                c_Body_y[1044] = n_Body_y[1044];
                c_Body_x[1045] = n_Body_x[1045];
                c_Body_y[1045] = n_Body_y[1045];
                c_Body_x[1046] = n_Body_x[1046];
                c_Body_y[1046] = n_Body_y[1046];
                c_Body_x[1047] = n_Body_x[1047];
                c_Body_y[1047] = n_Body_y[1047];
                c_Body_x[1048] = n_Body_x[1048];
                c_Body_y[1048] = n_Body_y[1048];
                c_Body_x[1049] = n_Body_x[1049];
                c_Body_y[1049] = n_Body_y[1049];
                c_Body_x[1050] = n_Body_x[1050];
                c_Body_y[1050] = n_Body_y[1050];
                c_Body_x[1051] = n_Body_x[1051];
                c_Body_y[1051] = n_Body_y[1051];
                c_Body_x[1052] = n_Body_x[1052];
                c_Body_y[1052] = n_Body_y[1052];
                c_Body_x[1053] = n_Body_x[1053];
                c_Body_y[1053] = n_Body_y[1053];
                c_Body_x[1054] = n_Body_x[1054];
                c_Body_y[1054] = n_Body_y[1054];
                c_Body_x[1055] = n_Body_x[1055];
                c_Body_y[1055] = n_Body_y[1055];
                c_Body_x[1056] = n_Body_x[1056];
                c_Body_y[1056] = n_Body_y[1056];
                c_Body_x[1057] = n_Body_x[1057];
                c_Body_y[1057] = n_Body_y[1057];
                c_Body_x[1058] = n_Body_x[1058];
                c_Body_y[1058] = n_Body_y[1058];
                c_Body_x[1059] = n_Body_x[1059];
                c_Body_y[1059] = n_Body_y[1059];
                c_Body_x[1060] = n_Body_x[1060];
                c_Body_y[1060] = n_Body_y[1060];
                c_Body_x[1061] = n_Body_x[1061];
                c_Body_y[1061] = n_Body_y[1061];
                c_Body_x[1062] = n_Body_x[1062];
                c_Body_y[1062] = n_Body_y[1062];
                c_Body_x[1063] = n_Body_x[1063];
                c_Body_y[1063] = n_Body_y[1063];
                c_Body_x[1064] = n_Body_x[1064];
                c_Body_y[1064] = n_Body_y[1064];
                c_Body_x[1065] = n_Body_x[1065];
                c_Body_y[1065] = n_Body_y[1065];
                c_Body_x[1066] = n_Body_x[1066];
                c_Body_y[1066] = n_Body_y[1066];
                c_Body_x[1067] = n_Body_x[1067];
                c_Body_y[1067] = n_Body_y[1067];
                c_Body_x[1068] = n_Body_x[1068];
                c_Body_y[1068] = n_Body_y[1068];
                c_Body_x[1069] = n_Body_x[1069];
                c_Body_y[1069] = n_Body_y[1069];
                c_Body_x[1070] = n_Body_x[1070];
                c_Body_y[1070] = n_Body_y[1070];
                c_Body_x[1071] = n_Body_x[1071];
                c_Body_y[1071] = n_Body_y[1071];
                c_Body_x[1072] = n_Body_x[1072];
                c_Body_y[1072] = n_Body_y[1072];
                c_Body_x[1073] = n_Body_x[1073];
                c_Body_y[1073] = n_Body_y[1073];
                c_Body_x[1074] = n_Body_x[1074];
                c_Body_y[1074] = n_Body_y[1074];
                c_Body_x[1075] = n_Body_x[1075];
                c_Body_y[1075] = n_Body_y[1075];
                c_Body_x[1076] = n_Body_x[1076];
                c_Body_y[1076] = n_Body_y[1076];
                c_Body_x[1077] = n_Body_x[1077];
                c_Body_y[1077] = n_Body_y[1077];
                c_Body_x[1078] = n_Body_x[1078];
                c_Body_y[1078] = n_Body_y[1078];
                c_Body_x[1079] = n_Body_x[1079];
                c_Body_y[1079] = n_Body_y[1079];
                c_Body_x[1080] = n_Body_x[1080];
                c_Body_y[1080] = n_Body_y[1080];
                c_Body_x[1081] = n_Body_x[1081];
                c_Body_y[1081] = n_Body_y[1081];
                c_Body_x[1082] = n_Body_x[1082];
                c_Body_y[1082] = n_Body_y[1082];
                c_Body_x[1083] = n_Body_x[1083];
                c_Body_y[1083] = n_Body_y[1083];
                c_Body_x[1084] = n_Body_x[1084];
                c_Body_y[1084] = n_Body_y[1084];
                c_Body_x[1085] = n_Body_x[1085];
                c_Body_y[1085] = n_Body_y[1085];
                c_Body_x[1086] = n_Body_x[1086];
                c_Body_y[1086] = n_Body_y[1086];
                c_Body_x[1087] = n_Body_x[1087];
                c_Body_y[1087] = n_Body_y[1087];
                c_Body_x[1088] = n_Body_x[1088];
                c_Body_y[1088] = n_Body_y[1088];
                c_Body_x[1089] = n_Body_x[1089];
                c_Body_y[1089] = n_Body_y[1089];
                c_Body_x[1090] = n_Body_x[1090];
                c_Body_y[1090] = n_Body_y[1090];
                c_Body_x[1091] = n_Body_x[1091];
                c_Body_y[1091] = n_Body_y[1091];
                c_Body_x[1092] = n_Body_x[1092];
                c_Body_y[1092] = n_Body_y[1092];
                c_Body_x[1093] = n_Body_x[1093];
                c_Body_y[1093] = n_Body_y[1093];
                c_Body_x[1094] = n_Body_x[1094];
                c_Body_y[1094] = n_Body_y[1094];
                c_Body_x[1095] = n_Body_x[1095];
                c_Body_y[1095] = n_Body_y[1095];
                c_Body_x[1096] = n_Body_x[1096];
                c_Body_y[1096] = n_Body_y[1096];
                c_Body_x[1097] = n_Body_x[1097];
                c_Body_y[1097] = n_Body_y[1097];
                c_Body_x[1098] = n_Body_x[1098];
                c_Body_y[1098] = n_Body_y[1098];
                c_Body_x[1099] = n_Body_x[1099];
                c_Body_y[1099] = n_Body_y[1099];
                c_Body_x[1100] = n_Body_x[1100];
                c_Body_y[1100] = n_Body_y[1100];
                c_Body_x[1101] = n_Body_x[1101];
                c_Body_y[1101] = n_Body_y[1101];
                c_Body_x[1102] = n_Body_x[1102];
                c_Body_y[1102] = n_Body_y[1102];
                c_Body_x[1103] = n_Body_x[1103];
                c_Body_y[1103] = n_Body_y[1103];
                c_Body_x[1104] = n_Body_x[1104];
                c_Body_y[1104] = n_Body_y[1104];
                c_Body_x[1105] = n_Body_x[1105];
                c_Body_y[1105] = n_Body_y[1105];
                c_Body_x[1106] = n_Body_x[1106];
                c_Body_y[1106] = n_Body_y[1106];
                c_Body_x[1107] = n_Body_x[1107];
                c_Body_y[1107] = n_Body_y[1107];
                c_Body_x[1108] = n_Body_x[1108];
                c_Body_y[1108] = n_Body_y[1108];
                c_Body_x[1109] = n_Body_x[1109];
                c_Body_y[1109] = n_Body_y[1109];
                c_Body_x[1110] = n_Body_x[1110];
                c_Body_y[1110] = n_Body_y[1110];
                c_Body_x[1111] = n_Body_x[1111];
                c_Body_y[1111] = n_Body_y[1111];
                c_Body_x[1112] = n_Body_x[1112];
                c_Body_y[1112] = n_Body_y[1112];
                c_Body_x[1113] = n_Body_x[1113];
                c_Body_y[1113] = n_Body_y[1113];
                c_Body_x[1114] = n_Body_x[1114];
                c_Body_y[1114] = n_Body_y[1114];
                c_Body_x[1115] = n_Body_x[1115];
                c_Body_y[1115] = n_Body_y[1115];
                c_Body_x[1116] = n_Body_x[1116];
                c_Body_y[1116] = n_Body_y[1116];
                c_Body_x[1117] = n_Body_x[1117];
                c_Body_y[1117] = n_Body_y[1117];
                c_Body_x[1118] = n_Body_x[1118];
                c_Body_y[1118] = n_Body_y[1118];
                c_Body_x[1119] = n_Body_x[1119];
                c_Body_y[1119] = n_Body_y[1119];
                c_Body_x[1120] = n_Body_x[1120];
                c_Body_y[1120] = n_Body_y[1120];
                c_Body_x[1121] = n_Body_x[1121];
                c_Body_y[1121] = n_Body_y[1121];
                c_Body_x[1122] = n_Body_x[1122];
                c_Body_y[1122] = n_Body_y[1122];
                c_Body_x[1123] = n_Body_x[1123];
                c_Body_y[1123] = n_Body_y[1123];
                c_Body_x[1124] = n_Body_x[1124];
                c_Body_y[1124] = n_Body_y[1124];
                c_Body_x[1125] = n_Body_x[1125];
                c_Body_y[1125] = n_Body_y[1125];
                c_Body_x[1126] = n_Body_x[1126];
                c_Body_y[1126] = n_Body_y[1126];
                c_Body_x[1127] = n_Body_x[1127];
                c_Body_y[1127] = n_Body_y[1127];
                c_Body_x[1128] = n_Body_x[1128];
                c_Body_y[1128] = n_Body_y[1128];
                c_Body_x[1129] = n_Body_x[1129];
                c_Body_y[1129] = n_Body_y[1129];
                c_Body_x[1130] = n_Body_x[1130];
                c_Body_y[1130] = n_Body_y[1130];
                c_Body_x[1131] = n_Body_x[1131];
                c_Body_y[1131] = n_Body_y[1131];
                c_Body_x[1132] = n_Body_x[1132];
                c_Body_y[1132] = n_Body_y[1132];
                c_Body_x[1133] = n_Body_x[1133];
                c_Body_y[1133] = n_Body_y[1133];
                c_Body_x[1134] = n_Body_x[1134];
                c_Body_y[1134] = n_Body_y[1134];
                c_Body_x[1135] = n_Body_x[1135];
                c_Body_y[1135] = n_Body_y[1135];
                c_Body_x[1136] = n_Body_x[1136];
                c_Body_y[1136] = n_Body_y[1136];
                c_Body_x[1137] = n_Body_x[1137];
                c_Body_y[1137] = n_Body_y[1137];
                c_Body_x[1138] = n_Body_x[1138];
                c_Body_y[1138] = n_Body_y[1138];
                c_Body_x[1139] = n_Body_x[1139];
                c_Body_y[1139] = n_Body_y[1139];
                c_Body_x[1140] = n_Body_x[1140];
                c_Body_y[1140] = n_Body_y[1140];
                c_Body_x[1141] = n_Body_x[1141];
                c_Body_y[1141] = n_Body_y[1141];
                c_Body_x[1142] = n_Body_x[1142];
                c_Body_y[1142] = n_Body_y[1142];
                c_Body_x[1143] = n_Body_x[1143];
                c_Body_y[1143] = n_Body_y[1143];
                c_Body_x[1144] = n_Body_x[1144];
                c_Body_y[1144] = n_Body_y[1144];
                c_Body_x[1145] = n_Body_x[1145];
                c_Body_y[1145] = n_Body_y[1145];
                c_Body_x[1146] = n_Body_x[1146];
                c_Body_y[1146] = n_Body_y[1146];
                c_Body_x[1147] = n_Body_x[1147];
                c_Body_y[1147] = n_Body_y[1147];
                c_Body_x[1148] = n_Body_x[1148];
                c_Body_y[1148] = n_Body_y[1148];
                c_Body_x[1149] = n_Body_x[1149];
                c_Body_y[1149] = n_Body_y[1149];
                c_Body_x[1150] = n_Body_x[1150];
                c_Body_y[1150] = n_Body_y[1150];
                c_Body_x[1151] = n_Body_x[1151];
                c_Body_y[1151] = n_Body_y[1151];
                c_Body_x[1152] = n_Body_x[1152];
                c_Body_y[1152] = n_Body_y[1152];
                c_Body_x[1153] = n_Body_x[1153];
                c_Body_y[1153] = n_Body_y[1153];
                c_Body_x[1154] = n_Body_x[1154];
                c_Body_y[1154] = n_Body_y[1154];
                c_Body_x[1155] = n_Body_x[1155];
                c_Body_y[1155] = n_Body_y[1155];
                c_Body_x[1156] = n_Body_x[1156];
                c_Body_y[1156] = n_Body_y[1156];
                c_Body_x[1157] = n_Body_x[1157];
                c_Body_y[1157] = n_Body_y[1157];
                c_Body_x[1158] = n_Body_x[1158];
                c_Body_y[1158] = n_Body_y[1158];
                c_Body_x[1159] = n_Body_x[1159];
                c_Body_y[1159] = n_Body_y[1159];
                c_Body_x[1160] = n_Body_x[1160];
                c_Body_y[1160] = n_Body_y[1160];
                c_Body_x[1161] = n_Body_x[1161];
                c_Body_y[1161] = n_Body_y[1161];
                c_Body_x[1162] = n_Body_x[1162];
                c_Body_y[1162] = n_Body_y[1162];
                c_Body_x[1163] = n_Body_x[1163];
                c_Body_y[1163] = n_Body_y[1163];
                c_Body_x[1164] = n_Body_x[1164];
                c_Body_y[1164] = n_Body_y[1164];
                c_Body_x[1165] = n_Body_x[1165];
                c_Body_y[1165] = n_Body_y[1165];
                c_Body_x[1166] = n_Body_x[1166];
                c_Body_y[1166] = n_Body_y[1166];
                c_Body_x[1167] = n_Body_x[1167];
                c_Body_y[1167] = n_Body_y[1167];
                c_Body_x[1168] = n_Body_x[1168];
                c_Body_y[1168] = n_Body_y[1168];
                c_Body_x[1169] = n_Body_x[1169];
                c_Body_y[1169] = n_Body_y[1169];
                c_Body_x[1170] = n_Body_x[1170];
                c_Body_y[1170] = n_Body_y[1170];
                c_Body_x[1171] = n_Body_x[1171];
                c_Body_y[1171] = n_Body_y[1171];
                c_Body_x[1172] = n_Body_x[1172];
                c_Body_y[1172] = n_Body_y[1172];
                c_Body_x[1173] = n_Body_x[1173];
                c_Body_y[1173] = n_Body_y[1173];
                c_Body_x[1174] = n_Body_x[1174];
                c_Body_y[1174] = n_Body_y[1174];
                c_Body_x[1175] = n_Body_x[1175];
                c_Body_y[1175] = n_Body_y[1175];
                c_Body_x[1176] = n_Body_x[1176];
                c_Body_y[1176] = n_Body_y[1176];
                c_Body_x[1177] = n_Body_x[1177];
                c_Body_y[1177] = n_Body_y[1177];
                c_Body_x[1178] = n_Body_x[1178];
                c_Body_y[1178] = n_Body_y[1178];
                c_Body_x[1179] = n_Body_x[1179];
                c_Body_y[1179] = n_Body_y[1179];
                c_Body_x[1180] = n_Body_x[1180];
                c_Body_y[1180] = n_Body_y[1180];
                c_Body_x[1181] = n_Body_x[1181];
                c_Body_y[1181] = n_Body_y[1181];
                c_Body_x[1182] = n_Body_x[1182];
                c_Body_y[1182] = n_Body_y[1182];
                c_Body_x[1183] = n_Body_x[1183];
                c_Body_y[1183] = n_Body_y[1183];
                c_Body_x[1184] = n_Body_x[1184];
                c_Body_y[1184] = n_Body_y[1184];
                c_Body_x[1185] = n_Body_x[1185];
                c_Body_y[1185] = n_Body_y[1185];
                c_Body_x[1186] = n_Body_x[1186];
                c_Body_y[1186] = n_Body_y[1186];
                c_Body_x[1187] = n_Body_x[1187];
                c_Body_y[1187] = n_Body_y[1187];
                c_Body_x[1188] = n_Body_x[1188];
                c_Body_y[1188] = n_Body_y[1188];
                c_Body_x[1189] = n_Body_x[1189];
                c_Body_y[1189] = n_Body_y[1189];
                c_Body_x[1190] = n_Body_x[1190];
                c_Body_y[1190] = n_Body_y[1190];
                c_Body_x[1191] = n_Body_x[1191];
                c_Body_y[1191] = n_Body_y[1191];
                c_Body_x[1192] = n_Body_x[1192];
                c_Body_y[1192] = n_Body_y[1192];
                c_Body_x[1193] = n_Body_x[1193];
                c_Body_y[1193] = n_Body_y[1193];
                c_Body_x[1194] = n_Body_x[1194];
                c_Body_y[1194] = n_Body_y[1194];
                c_Body_x[1195] = n_Body_x[1195];
                c_Body_y[1195] = n_Body_y[1195];
                c_Body_x[1196] = n_Body_x[1196];
                c_Body_y[1196] = n_Body_y[1196];
                c_Body_x[1197] = n_Body_x[1197];
                c_Body_y[1197] = n_Body_y[1197];
                c_Body_x[1198] = n_Body_x[1198];
                c_Body_y[1198] = n_Body_y[1198];
                c_Body_x[1199] = n_Body_x[1199];
                c_Body_y[1199] = n_Body_y[1199];
                c_Body_x[1200] = n_Body_x[1200];
                c_Body_y[1200] = n_Body_y[1200];
                c_Body_x[1201] = n_Body_x[1201];
                c_Body_y[1201] = n_Body_y[1201];
                c_Body_x[1202] = n_Body_x[1202];
                c_Body_y[1202] = n_Body_y[1202];
                c_Body_x[1203] = n_Body_x[1203];
                c_Body_y[1203] = n_Body_y[1203];
                c_Body_x[1204] = n_Body_x[1204];
                c_Body_y[1204] = n_Body_y[1204];
                c_Body_x[1205] = n_Body_x[1205];
                c_Body_y[1205] = n_Body_y[1205];
                c_Body_x[1206] = n_Body_x[1206];
                c_Body_y[1206] = n_Body_y[1206];
                c_Body_x[1207] = n_Body_x[1207];
                c_Body_y[1207] = n_Body_y[1207];
                c_Body_x[1208] = n_Body_x[1208];
                c_Body_y[1208] = n_Body_y[1208];
                c_Body_x[1209] = n_Body_x[1209];
                c_Body_y[1209] = n_Body_y[1209];
                c_Body_x[1210] = n_Body_x[1210];
                c_Body_y[1210] = n_Body_y[1210];
                c_Body_x[1211] = n_Body_x[1211];
                c_Body_y[1211] = n_Body_y[1211];
                c_Body_x[1212] = n_Body_x[1212];
                c_Body_y[1212] = n_Body_y[1212];
                c_Body_x[1213] = n_Body_x[1213];
                c_Body_y[1213] = n_Body_y[1213];
                c_Body_x[1214] = n_Body_x[1214];
                c_Body_y[1214] = n_Body_y[1214];
                c_Body_x[1215] = n_Body_x[1215];
                c_Body_y[1215] = n_Body_y[1215];
                c_Body_x[1216] = n_Body_x[1216];
                c_Body_y[1216] = n_Body_y[1216];
                c_Body_x[1217] = n_Body_x[1217];
                c_Body_y[1217] = n_Body_y[1217];
                c_Body_x[1218] = n_Body_x[1218];
                c_Body_y[1218] = n_Body_y[1218];
                c_Body_x[1219] = n_Body_x[1219];
                c_Body_y[1219] = n_Body_y[1219];
                c_Body_x[1220] = n_Body_x[1220];
                c_Body_y[1220] = n_Body_y[1220];
                c_Body_x[1221] = n_Body_x[1221];
                c_Body_y[1221] = n_Body_y[1221];
                c_Body_x[1222] = n_Body_x[1222];
                c_Body_y[1222] = n_Body_y[1222];
                c_Body_x[1223] = n_Body_x[1223];
                c_Body_y[1223] = n_Body_y[1223];
                c_Body_x[1224] = n_Body_x[1224];
                c_Body_y[1224] = n_Body_y[1224];
                c_Body_x[1225] = n_Body_x[1225];
                c_Body_y[1225] = n_Body_y[1225];
                c_Body_x[1226] = n_Body_x[1226];
                c_Body_y[1226] = n_Body_y[1226];
                c_Body_x[1227] = n_Body_x[1227];
                c_Body_y[1227] = n_Body_y[1227];
                c_Body_x[1228] = n_Body_x[1228];
                c_Body_y[1228] = n_Body_y[1228];
                c_Body_x[1229] = n_Body_x[1229];
                c_Body_y[1229] = n_Body_y[1229];
                c_Body_x[1230] = n_Body_x[1230];
                c_Body_y[1230] = n_Body_y[1230];
                c_Body_x[1231] = n_Body_x[1231];
                c_Body_y[1231] = n_Body_y[1231];
                c_Body_x[1232] = n_Body_x[1232];
                c_Body_y[1232] = n_Body_y[1232];
                c_Body_x[1233] = n_Body_x[1233];
                c_Body_y[1233] = n_Body_y[1233];
                c_Body_x[1234] = n_Body_x[1234];
                c_Body_y[1234] = n_Body_y[1234];
                c_Body_x[1235] = n_Body_x[1235];
                c_Body_y[1235] = n_Body_y[1235];
                c_Body_x[1236] = n_Body_x[1236];
                c_Body_y[1236] = n_Body_y[1236];
                c_Body_x[1237] = n_Body_x[1237];
                c_Body_y[1237] = n_Body_y[1237];
                c_Body_x[1238] = n_Body_x[1238];
                c_Body_y[1238] = n_Body_y[1238];
                c_Body_x[1239] = n_Body_x[1239];
                c_Body_y[1239] = n_Body_y[1239];
                c_Body_x[1240] = n_Body_x[1240];
                c_Body_y[1240] = n_Body_y[1240];
                c_Body_x[1241] = n_Body_x[1241];
                c_Body_y[1241] = n_Body_y[1241];
                c_Body_x[1242] = n_Body_x[1242];
                c_Body_y[1242] = n_Body_y[1242];
                c_Body_x[1243] = n_Body_x[1243];
                c_Body_y[1243] = n_Body_y[1243];
                c_Body_x[1244] = n_Body_x[1244];
                c_Body_y[1244] = n_Body_y[1244];
                c_Body_x[1245] = n_Body_x[1245];
                c_Body_y[1245] = n_Body_y[1245];
                c_Body_x[1246] = n_Body_x[1246];
                c_Body_y[1246] = n_Body_y[1246];
                c_Body_x[1247] = n_Body_x[1247];
                c_Body_y[1247] = n_Body_y[1247];
                c_Body_x[1248] = n_Body_x[1248];
                c_Body_y[1248] = n_Body_y[1248];
                c_Body_x[1249] = n_Body_x[1249];
                c_Body_y[1249] = n_Body_y[1249];
                c_Body_x[1250] = n_Body_x[1250];
                c_Body_y[1250] = n_Body_y[1250];
                c_Body_x[1251] = n_Body_x[1251];
                c_Body_y[1251] = n_Body_y[1251];
                c_Body_x[1252] = n_Body_x[1252];
                c_Body_y[1252] = n_Body_y[1252];
                c_Body_x[1253] = n_Body_x[1253];
                c_Body_y[1253] = n_Body_y[1253];
                c_Body_x[1254] = n_Body_x[1254];
                c_Body_y[1254] = n_Body_y[1254];
                c_Body_x[1255] = n_Body_x[1255];
                c_Body_y[1255] = n_Body_y[1255];
                c_Body_x[1256] = n_Body_x[1256];
                c_Body_y[1256] = n_Body_y[1256];
                c_Body_x[1257] = n_Body_x[1257];
                c_Body_y[1257] = n_Body_y[1257];
                c_Body_x[1258] = n_Body_x[1258];
                c_Body_y[1258] = n_Body_y[1258];
                c_Body_x[1259] = n_Body_x[1259];
                c_Body_y[1259] = n_Body_y[1259];
                c_Body_x[1260] = n_Body_x[1260];
                c_Body_y[1260] = n_Body_y[1260];
                c_Body_x[1261] = n_Body_x[1261];
                c_Body_y[1261] = n_Body_y[1261];
                c_Body_x[1262] = n_Body_x[1262];
                c_Body_y[1262] = n_Body_y[1262];
                c_Body_x[1263] = n_Body_x[1263];
                c_Body_y[1263] = n_Body_y[1263];
                c_Body_x[1264] = n_Body_x[1264];
                c_Body_y[1264] = n_Body_y[1264];
                c_Body_x[1265] = n_Body_x[1265];
                c_Body_y[1265] = n_Body_y[1265];
                c_Body_x[1266] = n_Body_x[1266];
                c_Body_y[1266] = n_Body_y[1266];
                c_Body_x[1267] = n_Body_x[1267];
                c_Body_y[1267] = n_Body_y[1267];
                c_Body_x[1268] = n_Body_x[1268];
                c_Body_y[1268] = n_Body_y[1268];
                c_Body_x[1269] = n_Body_x[1269];
                c_Body_y[1269] = n_Body_y[1269];
                c_Body_x[1270] = n_Body_x[1270];
                c_Body_y[1270] = n_Body_y[1270];
                c_Body_x[1271] = n_Body_x[1271];
                c_Body_y[1271] = n_Body_y[1271];
                c_Body_x[1272] = n_Body_x[1272];
                c_Body_y[1272] = n_Body_y[1272];
                c_Body_x[1273] = n_Body_x[1273];
                c_Body_y[1273] = n_Body_y[1273];
                c_Body_x[1274] = n_Body_x[1274];
                c_Body_y[1274] = n_Body_y[1274];
                c_Body_x[1275] = n_Body_x[1275];
                c_Body_y[1275] = n_Body_y[1275];
                c_Body_x[1276] = n_Body_x[1276];
                c_Body_y[1276] = n_Body_y[1276];
                c_Body_x[1277] = n_Body_x[1277];
                c_Body_y[1277] = n_Body_y[1277];
                c_Body_x[1278] = n_Body_x[1278];
                c_Body_y[1278] = n_Body_y[1278];
                c_Body_x[1279] = n_Body_x[1279];
                c_Body_y[1279] = n_Body_y[1279];
                c_Body_x[1280] = n_Body_x[1280];
                c_Body_y[1280] = n_Body_y[1280];
                c_Body_x[1281] = n_Body_x[1281];
                c_Body_y[1281] = n_Body_y[1281];
                c_Body_x[1282] = n_Body_x[1282];
                c_Body_y[1282] = n_Body_y[1282];
                c_Body_x[1283] = n_Body_x[1283];
                c_Body_y[1283] = n_Body_y[1283];
                c_Body_x[1284] = n_Body_x[1284];
                c_Body_y[1284] = n_Body_y[1284];
                c_Body_x[1285] = n_Body_x[1285];
                c_Body_y[1285] = n_Body_y[1285];
                c_Body_x[1286] = n_Body_x[1286];
                c_Body_y[1286] = n_Body_y[1286];
                c_Body_x[1287] = n_Body_x[1287];
                c_Body_y[1287] = n_Body_y[1287];
                c_Body_x[1288] = n_Body_x[1288];
                c_Body_y[1288] = n_Body_y[1288];
                c_Body_x[1289] = n_Body_x[1289];
                c_Body_y[1289] = n_Body_y[1289];
                c_Body_x[1290] = n_Body_x[1290];
                c_Body_y[1290] = n_Body_y[1290];
                c_Body_x[1291] = n_Body_x[1291];
                c_Body_y[1291] = n_Body_y[1291];
                c_Body_x[1292] = n_Body_x[1292];
                c_Body_y[1292] = n_Body_y[1292];
                c_Body_x[1293] = n_Body_x[1293];
                c_Body_y[1293] = n_Body_y[1293];
                c_Body_x[1294] = n_Body_x[1294];
                c_Body_y[1294] = n_Body_y[1294];
                c_Body_x[1295] = n_Body_x[1295];
                c_Body_y[1295] = n_Body_y[1295];
                c_Body_x[1296] = n_Body_x[1296];
                c_Body_y[1296] = n_Body_y[1296];
                c_Body_x[1297] = n_Body_x[1297];
                c_Body_y[1297] = n_Body_y[1297];
                c_Body_x[1298] = n_Body_x[1298];
                c_Body_y[1298] = n_Body_y[1298];
                c_Body_x[1299] = n_Body_x[1299];
                c_Body_y[1299] = n_Body_y[1299];
                c_Body_x[1300] = n_Body_x[1300];
                c_Body_y[1300] = n_Body_y[1300];
                c_Body_x[1301] = n_Body_x[1301];
                c_Body_y[1301] = n_Body_y[1301];
                c_Body_x[1302] = n_Body_x[1302];
                c_Body_y[1302] = n_Body_y[1302];
                c_Body_x[1303] = n_Body_x[1303];
                c_Body_y[1303] = n_Body_y[1303];
                c_Body_x[1304] = n_Body_x[1304];
                c_Body_y[1304] = n_Body_y[1304];
                c_Body_x[1305] = n_Body_x[1305];
                c_Body_y[1305] = n_Body_y[1305];
                c_Body_x[1306] = n_Body_x[1306];
                c_Body_y[1306] = n_Body_y[1306];
                c_Body_x[1307] = n_Body_x[1307];
                c_Body_y[1307] = n_Body_y[1307];
                c_Body_x[1308] = n_Body_x[1308];
                c_Body_y[1308] = n_Body_y[1308];
                c_Body_x[1309] = n_Body_x[1309];
                c_Body_y[1309] = n_Body_y[1309];
                c_Body_x[1310] = n_Body_x[1310];
                c_Body_y[1310] = n_Body_y[1310];
                c_Body_x[1311] = n_Body_x[1311];
                c_Body_y[1311] = n_Body_y[1311];
                c_Body_x[1312] = n_Body_x[1312];
                c_Body_y[1312] = n_Body_y[1312];
                c_Body_x[1313] = n_Body_x[1313];
                c_Body_y[1313] = n_Body_y[1313];
                c_Body_x[1314] = n_Body_x[1314];
                c_Body_y[1314] = n_Body_y[1314];
                c_Body_x[1315] = n_Body_x[1315];
                c_Body_y[1315] = n_Body_y[1315];
                c_Body_x[1316] = n_Body_x[1316];
                c_Body_y[1316] = n_Body_y[1316];
                c_Body_x[1317] = n_Body_x[1317];
                c_Body_y[1317] = n_Body_y[1317];
                c_Body_x[1318] = n_Body_x[1318];
                c_Body_y[1318] = n_Body_y[1318];
                c_Body_x[1319] = n_Body_x[1319];
                c_Body_y[1319] = n_Body_y[1319];
                c_Body_x[1320] = n_Body_x[1320];
                c_Body_y[1320] = n_Body_y[1320];
                c_Body_x[1321] = n_Body_x[1321];
                c_Body_y[1321] = n_Body_y[1321];
                c_Body_x[1322] = n_Body_x[1322];
                c_Body_y[1322] = n_Body_y[1322];
                c_Body_x[1323] = n_Body_x[1323];
                c_Body_y[1323] = n_Body_y[1323];
                c_Body_x[1324] = n_Body_x[1324];
                c_Body_y[1324] = n_Body_y[1324];
                c_Body_x[1325] = n_Body_x[1325];
                c_Body_y[1325] = n_Body_y[1325];
                c_Body_x[1326] = n_Body_x[1326];
                c_Body_y[1326] = n_Body_y[1326];
                c_Body_x[1327] = n_Body_x[1327];
                c_Body_y[1327] = n_Body_y[1327];
                c_Body_x[1328] = n_Body_x[1328];
                c_Body_y[1328] = n_Body_y[1328];
                c_Body_x[1329] = n_Body_x[1329];
                c_Body_y[1329] = n_Body_y[1329];
                c_Body_x[1330] = n_Body_x[1330];
                c_Body_y[1330] = n_Body_y[1330];
                c_Body_x[1331] = n_Body_x[1331];
                c_Body_y[1331] = n_Body_y[1331];
                c_Body_x[1332] = n_Body_x[1332];
                c_Body_y[1332] = n_Body_y[1332];
                c_Body_x[1333] = n_Body_x[1333];
                c_Body_y[1333] = n_Body_y[1333];
                c_Body_x[1334] = n_Body_x[1334];
                c_Body_y[1334] = n_Body_y[1334];
                c_Body_x[1335] = n_Body_x[1335];
                c_Body_y[1335] = n_Body_y[1335];
                c_Body_x[1336] = n_Body_x[1336];
                c_Body_y[1336] = n_Body_y[1336];
                c_Body_x[1337] = n_Body_x[1337];
                c_Body_y[1337] = n_Body_y[1337];
                c_Body_x[1338] = n_Body_x[1338];
                c_Body_y[1338] = n_Body_y[1338];
                c_Body_x[1339] = n_Body_x[1339];
                c_Body_y[1339] = n_Body_y[1339];
                c_Body_x[1340] = n_Body_x[1340];
                c_Body_y[1340] = n_Body_y[1340];
                c_Body_x[1341] = n_Body_x[1341];
                c_Body_y[1341] = n_Body_y[1341];
                c_Body_x[1342] = n_Body_x[1342];
                c_Body_y[1342] = n_Body_y[1342];
                c_Body_x[1343] = n_Body_x[1343];
                c_Body_y[1343] = n_Body_y[1343];
                c_Body_x[1344] = n_Body_x[1344];
                c_Body_y[1344] = n_Body_y[1344];
                c_Body_x[1345] = n_Body_x[1345];
                c_Body_y[1345] = n_Body_y[1345];
                c_Body_x[1346] = n_Body_x[1346];
                c_Body_y[1346] = n_Body_y[1346];
                c_Body_x[1347] = n_Body_x[1347];
                c_Body_y[1347] = n_Body_y[1347];
                c_Body_x[1348] = n_Body_x[1348];
                c_Body_y[1348] = n_Body_y[1348];
                c_Body_x[1349] = n_Body_x[1349];
                c_Body_y[1349] = n_Body_y[1349];
                c_Body_x[1350] = n_Body_x[1350];
                c_Body_y[1350] = n_Body_y[1350];
                c_Body_x[1351] = n_Body_x[1351];
                c_Body_y[1351] = n_Body_y[1351];
                c_Body_x[1352] = n_Body_x[1352];
                c_Body_y[1352] = n_Body_y[1352];
                c_Body_x[1353] = n_Body_x[1353];
                c_Body_y[1353] = n_Body_y[1353];
                c_Body_x[1354] = n_Body_x[1354];
                c_Body_y[1354] = n_Body_y[1354];
                c_Body_x[1355] = n_Body_x[1355];
                c_Body_y[1355] = n_Body_y[1355];
                c_Body_x[1356] = n_Body_x[1356];
                c_Body_y[1356] = n_Body_y[1356];
                c_Body_x[1357] = n_Body_x[1357];
                c_Body_y[1357] = n_Body_y[1357];
                c_Body_x[1358] = n_Body_x[1358];
                c_Body_y[1358] = n_Body_y[1358];
                c_Body_x[1359] = n_Body_x[1359];
                c_Body_y[1359] = n_Body_y[1359];
                c_Body_x[1360] = n_Body_x[1360];
                c_Body_y[1360] = n_Body_y[1360];
                c_Body_x[1361] = n_Body_x[1361];
                c_Body_y[1361] = n_Body_y[1361];
                c_Body_x[1362] = n_Body_x[1362];
                c_Body_y[1362] = n_Body_y[1362];
                c_Body_x[1363] = n_Body_x[1363];
                c_Body_y[1363] = n_Body_y[1363];
                c_Body_x[1364] = n_Body_x[1364];
                c_Body_y[1364] = n_Body_y[1364];
                c_Body_x[1365] = n_Body_x[1365];
                c_Body_y[1365] = n_Body_y[1365];
                c_Body_x[1366] = n_Body_x[1366];
                c_Body_y[1366] = n_Body_y[1366];
                c_Body_x[1367] = n_Body_x[1367];
                c_Body_y[1367] = n_Body_y[1367];
                c_Body_x[1368] = n_Body_x[1368];
                c_Body_y[1368] = n_Body_y[1368];
                c_Body_x[1369] = n_Body_x[1369];
                c_Body_y[1369] = n_Body_y[1369];
                c_Body_x[1370] = n_Body_x[1370];
                c_Body_y[1370] = n_Body_y[1370];
                c_Body_x[1371] = n_Body_x[1371];
                c_Body_y[1371] = n_Body_y[1371];
                c_Body_x[1372] = n_Body_x[1372];
                c_Body_y[1372] = n_Body_y[1372];
                c_Body_x[1373] = n_Body_x[1373];
                c_Body_y[1373] = n_Body_y[1373];
                c_Body_x[1374] = n_Body_x[1374];
                c_Body_y[1374] = n_Body_y[1374];
                c_Body_x[1375] = n_Body_x[1375];
                c_Body_y[1375] = n_Body_y[1375];
                c_Body_x[1376] = n_Body_x[1376];
                c_Body_y[1376] = n_Body_y[1376];
                c_Body_x[1377] = n_Body_x[1377];
                c_Body_y[1377] = n_Body_y[1377];
                c_Body_x[1378] = n_Body_x[1378];
                c_Body_y[1378] = n_Body_y[1378];
                c_Body_x[1379] = n_Body_x[1379];
                c_Body_y[1379] = n_Body_y[1379];
                c_Body_x[1380] = n_Body_x[1380];
                c_Body_y[1380] = n_Body_y[1380];
                c_Body_x[1381] = n_Body_x[1381];
                c_Body_y[1381] = n_Body_y[1381];
                c_Body_x[1382] = n_Body_x[1382];
                c_Body_y[1382] = n_Body_y[1382];
                c_Body_x[1383] = n_Body_x[1383];
                c_Body_y[1383] = n_Body_y[1383];
                c_Body_x[1384] = n_Body_x[1384];
                c_Body_y[1384] = n_Body_y[1384];
                c_Body_x[1385] = n_Body_x[1385];
                c_Body_y[1385] = n_Body_y[1385];
                c_Body_x[1386] = n_Body_x[1386];
                c_Body_y[1386] = n_Body_y[1386];
                c_Body_x[1387] = n_Body_x[1387];
                c_Body_y[1387] = n_Body_y[1387];
                c_Body_x[1388] = n_Body_x[1388];
                c_Body_y[1388] = n_Body_y[1388];
                c_Body_x[1389] = n_Body_x[1389];
                c_Body_y[1389] = n_Body_y[1389];
                c_Body_x[1390] = n_Body_x[1390];
                c_Body_y[1390] = n_Body_y[1390];
                c_Body_x[1391] = n_Body_x[1391];
                c_Body_y[1391] = n_Body_y[1391];
                c_Body_x[1392] = n_Body_x[1392];
                c_Body_y[1392] = n_Body_y[1392];
                c_Body_x[1393] = n_Body_x[1393];
                c_Body_y[1393] = n_Body_y[1393];
                c_Body_x[1394] = n_Body_x[1394];
                c_Body_y[1394] = n_Body_y[1394];
                c_Body_x[1395] = n_Body_x[1395];
                c_Body_y[1395] = n_Body_y[1395];
                c_Body_x[1396] = n_Body_x[1396];
                c_Body_y[1396] = n_Body_y[1396];
                c_Body_x[1397] = n_Body_x[1397];
                c_Body_y[1397] = n_Body_y[1397];
                c_Body_x[1398] = n_Body_x[1398];
                c_Body_y[1398] = n_Body_y[1398];
                c_Body_x[1399] = n_Body_x[1399];
                c_Body_y[1399] = n_Body_y[1399];
                c_Body_x[1400] = n_Body_x[1400];
                c_Body_y[1400] = n_Body_y[1400];
                c_Body_x[1401] = n_Body_x[1401];
                c_Body_y[1401] = n_Body_y[1401];
                c_Body_x[1402] = n_Body_x[1402];
                c_Body_y[1402] = n_Body_y[1402];
                c_Body_x[1403] = n_Body_x[1403];
                c_Body_y[1403] = n_Body_y[1403];
                c_Body_x[1404] = n_Body_x[1404];
                c_Body_y[1404] = n_Body_y[1404];
                c_Body_x[1405] = n_Body_x[1405];
                c_Body_y[1405] = n_Body_y[1405];
                c_Body_x[1406] = n_Body_x[1406];
                c_Body_y[1406] = n_Body_y[1406];
                c_Body_x[1407] = n_Body_x[1407];
                c_Body_y[1407] = n_Body_y[1407];
                c_Body_x[1408] = n_Body_x[1408];
                c_Body_y[1408] = n_Body_y[1408];
                c_Body_x[1409] = n_Body_x[1409];
                c_Body_y[1409] = n_Body_y[1409];
                c_Body_x[1410] = n_Body_x[1410];
                c_Body_y[1410] = n_Body_y[1410];
                c_Body_x[1411] = n_Body_x[1411];
                c_Body_y[1411] = n_Body_y[1411];
                c_Body_x[1412] = n_Body_x[1412];
                c_Body_y[1412] = n_Body_y[1412];
                c_Body_x[1413] = n_Body_x[1413];
                c_Body_y[1413] = n_Body_y[1413];
                c_Body_x[1414] = n_Body_x[1414];
                c_Body_y[1414] = n_Body_y[1414];
                c_Body_x[1415] = n_Body_x[1415];
                c_Body_y[1415] = n_Body_y[1415];
                c_Body_x[1416] = n_Body_x[1416];
                c_Body_y[1416] = n_Body_y[1416];
                c_Body_x[1417] = n_Body_x[1417];
                c_Body_y[1417] = n_Body_y[1417];
                c_Body_x[1418] = n_Body_x[1418];
                c_Body_y[1418] = n_Body_y[1418];
                c_Body_x[1419] = n_Body_x[1419];
                c_Body_y[1419] = n_Body_y[1419];
                c_Body_x[1420] = n_Body_x[1420];
                c_Body_y[1420] = n_Body_y[1420];
                c_Body_x[1421] = n_Body_x[1421];
                c_Body_y[1421] = n_Body_y[1421];
                c_Body_x[1422] = n_Body_x[1422];
                c_Body_y[1422] = n_Body_y[1422];
                c_Body_x[1423] = n_Body_x[1423];
                c_Body_y[1423] = n_Body_y[1423];
                c_Body_x[1424] = n_Body_x[1424];
                c_Body_y[1424] = n_Body_y[1424];
                c_Body_x[1425] = n_Body_x[1425];
                c_Body_y[1425] = n_Body_y[1425];
                c_Body_x[1426] = n_Body_x[1426];
                c_Body_y[1426] = n_Body_y[1426];
                c_Body_x[1427] = n_Body_x[1427];
                c_Body_y[1427] = n_Body_y[1427];
                c_Body_x[1428] = n_Body_x[1428];
                c_Body_y[1428] = n_Body_y[1428];
                c_Body_x[1429] = n_Body_x[1429];
                c_Body_y[1429] = n_Body_y[1429];
                c_Body_x[1430] = n_Body_x[1430];
                c_Body_y[1430] = n_Body_y[1430];
                c_Body_x[1431] = n_Body_x[1431];
                c_Body_y[1431] = n_Body_y[1431];
                c_Body_x[1432] = n_Body_x[1432];
                c_Body_y[1432] = n_Body_y[1432];
                c_Body_x[1433] = n_Body_x[1433];
                c_Body_y[1433] = n_Body_y[1433];
                c_Body_x[1434] = n_Body_x[1434];
                c_Body_y[1434] = n_Body_y[1434];
                c_Body_x[1435] = n_Body_x[1435];
                c_Body_y[1435] = n_Body_y[1435];
                c_Body_x[1436] = n_Body_x[1436];
                c_Body_y[1436] = n_Body_y[1436];
                c_Body_x[1437] = n_Body_x[1437];
                c_Body_y[1437] = n_Body_y[1437];
                c_Body_x[1438] = n_Body_x[1438];
                c_Body_y[1438] = n_Body_y[1438];
                c_Body_x[1439] = n_Body_x[1439];
                c_Body_y[1439] = n_Body_y[1439];
                c_Body_x[1440] = n_Body_x[1440];
                c_Body_y[1440] = n_Body_y[1440];
                c_Body_x[1441] = n_Body_x[1441];
                c_Body_y[1441] = n_Body_y[1441];
                c_Body_x[1442] = n_Body_x[1442];
                c_Body_y[1442] = n_Body_y[1442];
                c_Body_x[1443] = n_Body_x[1443];
                c_Body_y[1443] = n_Body_y[1443];
                c_Body_x[1444] = n_Body_x[1444];
                c_Body_y[1444] = n_Body_y[1444];
                c_Body_x[1445] = n_Body_x[1445];
                c_Body_y[1445] = n_Body_y[1445];
                c_Body_x[1446] = n_Body_x[1446];
                c_Body_y[1446] = n_Body_y[1446];
                c_Body_x[1447] = n_Body_x[1447];
                c_Body_y[1447] = n_Body_y[1447];
                c_Body_x[1448] = n_Body_x[1448];
                c_Body_y[1448] = n_Body_y[1448];
                c_Body_x[1449] = n_Body_x[1449];
                c_Body_y[1449] = n_Body_y[1449];
                c_Body_x[1450] = n_Body_x[1450];
                c_Body_y[1450] = n_Body_y[1450];
                c_Body_x[1451] = n_Body_x[1451];
                c_Body_y[1451] = n_Body_y[1451];
                c_Body_x[1452] = n_Body_x[1452];
                c_Body_y[1452] = n_Body_y[1452];
                c_Body_x[1453] = n_Body_x[1453];
                c_Body_y[1453] = n_Body_y[1453];
                c_Body_x[1454] = n_Body_x[1454];
                c_Body_y[1454] = n_Body_y[1454];
                c_Body_x[1455] = n_Body_x[1455];
                c_Body_y[1455] = n_Body_y[1455];
                c_Body_x[1456] = n_Body_x[1456];
                c_Body_y[1456] = n_Body_y[1456];
                c_Body_x[1457] = n_Body_x[1457];
                c_Body_y[1457] = n_Body_y[1457];
                c_Body_x[1458] = n_Body_x[1458];
                c_Body_y[1458] = n_Body_y[1458];
                c_Body_x[1459] = n_Body_x[1459];
                c_Body_y[1459] = n_Body_y[1459];
                c_Body_x[1460] = n_Body_x[1460];
                c_Body_y[1460] = n_Body_y[1460];
                c_Body_x[1461] = n_Body_x[1461];
                c_Body_y[1461] = n_Body_y[1461];
                c_Body_x[1462] = n_Body_x[1462];
                c_Body_y[1462] = n_Body_y[1462];
                c_Body_x[1463] = n_Body_x[1463];
                c_Body_y[1463] = n_Body_y[1463];
                c_Body_x[1464] = n_Body_x[1464];
                c_Body_y[1464] = n_Body_y[1464];
                c_Body_x[1465] = n_Body_x[1465];
                c_Body_y[1465] = n_Body_y[1465];
                c_Body_x[1466] = n_Body_x[1466];
                c_Body_y[1466] = n_Body_y[1466];
                c_Body_x[1467] = n_Body_x[1467];
                c_Body_y[1467] = n_Body_y[1467];
                c_Body_x[1468] = n_Body_x[1468];
                c_Body_y[1468] = n_Body_y[1468];
                c_Body_x[1469] = n_Body_x[1469];
                c_Body_y[1469] = n_Body_y[1469];
                c_Body_x[1470] = n_Body_x[1470];
                c_Body_y[1470] = n_Body_y[1470];
                c_Body_x[1471] = n_Body_x[1471];
                c_Body_y[1471] = n_Body_y[1471];
                c_Body_x[1472] = n_Body_x[1472];
                c_Body_y[1472] = n_Body_y[1472];
                c_Body_x[1473] = n_Body_x[1473];
                c_Body_y[1473] = n_Body_y[1473];
                c_Body_x[1474] = n_Body_x[1474];
                c_Body_y[1474] = n_Body_y[1474];
                c_Body_x[1475] = n_Body_x[1475];
                c_Body_y[1475] = n_Body_y[1475];
                c_Body_x[1476] = n_Body_x[1476];
                c_Body_y[1476] = n_Body_y[1476];
                c_Body_x[1477] = n_Body_x[1477];
                c_Body_y[1477] = n_Body_y[1477];
                c_Body_x[1478] = n_Body_x[1478];
                c_Body_y[1478] = n_Body_y[1478];
                c_Body_x[1479] = n_Body_x[1479];
                c_Body_y[1479] = n_Body_y[1479];
                c_Body_x[1480] = n_Body_x[1480];
                c_Body_y[1480] = n_Body_y[1480];
                c_Body_x[1481] = n_Body_x[1481];
                c_Body_y[1481] = n_Body_y[1481];
                c_Body_x[1482] = n_Body_x[1482];
                c_Body_y[1482] = n_Body_y[1482];
                c_Body_x[1483] = n_Body_x[1483];
                c_Body_y[1483] = n_Body_y[1483];
                c_Body_x[1484] = n_Body_x[1484];
                c_Body_y[1484] = n_Body_y[1484];
                c_Body_x[1485] = n_Body_x[1485];
                c_Body_y[1485] = n_Body_y[1485];
                c_Body_x[1486] = n_Body_x[1486];
                c_Body_y[1486] = n_Body_y[1486];
                c_Body_x[1487] = n_Body_x[1487];
                c_Body_y[1487] = n_Body_y[1487];
                c_Body_x[1488] = n_Body_x[1488];
                c_Body_y[1488] = n_Body_y[1488];
                c_Body_x[1489] = n_Body_x[1489];
                c_Body_y[1489] = n_Body_y[1489];
                c_Body_x[1490] = n_Body_x[1490];
                c_Body_y[1490] = n_Body_y[1490];
                c_Body_x[1491] = n_Body_x[1491];
                c_Body_y[1491] = n_Body_y[1491];
                c_Body_x[1492] = n_Body_x[1492];
                c_Body_y[1492] = n_Body_y[1492];
                c_Body_x[1493] = n_Body_x[1493];
                c_Body_y[1493] = n_Body_y[1493];
                c_Body_x[1494] = n_Body_x[1494];
                c_Body_y[1494] = n_Body_y[1494];
                c_Body_x[1495] = n_Body_x[1495];
                c_Body_y[1495] = n_Body_y[1495];
                c_Body_x[1496] = n_Body_x[1496];
                c_Body_y[1496] = n_Body_y[1496];
                c_Body_x[1497] = n_Body_x[1497];
                c_Body_y[1497] = n_Body_y[1497];
                c_Body_x[1498] = n_Body_x[1498];
                c_Body_y[1498] = n_Body_y[1498];
                c_Body_x[1499] = n_Body_x[1499];
                c_Body_y[1499] = n_Body_y[1499];
                c_Body_x[1500] = n_Body_x[1500];
                c_Body_y[1500] = n_Body_y[1500];
                c_Body_x[1501] = n_Body_x[1501];
                c_Body_y[1501] = n_Body_y[1501];
                c_Body_x[1502] = n_Body_x[1502];
                c_Body_y[1502] = n_Body_y[1502];
                c_Body_x[1503] = n_Body_x[1503];
                c_Body_y[1503] = n_Body_y[1503];
                c_Body_x[1504] = n_Body_x[1504];
                c_Body_y[1504] = n_Body_y[1504];
                c_Body_x[1505] = n_Body_x[1505];
                c_Body_y[1505] = n_Body_y[1505];
                c_Body_x[1506] = n_Body_x[1506];
                c_Body_y[1506] = n_Body_y[1506];
                c_Body_x[1507] = n_Body_x[1507];
                c_Body_y[1507] = n_Body_y[1507];
                c_Body_x[1508] = n_Body_x[1508];
                c_Body_y[1508] = n_Body_y[1508];
                c_Body_x[1509] = n_Body_x[1509];
                c_Body_y[1509] = n_Body_y[1509];
                c_Body_x[1510] = n_Body_x[1510];
                c_Body_y[1510] = n_Body_y[1510];
                c_Body_x[1511] = n_Body_x[1511];
                c_Body_y[1511] = n_Body_y[1511];
                c_Body_x[1512] = n_Body_x[1512];
                c_Body_y[1512] = n_Body_y[1512];
                c_Body_x[1513] = n_Body_x[1513];
                c_Body_y[1513] = n_Body_y[1513];
                c_Body_x[1514] = n_Body_x[1514];
                c_Body_y[1514] = n_Body_y[1514];
                c_Body_x[1515] = n_Body_x[1515];
                c_Body_y[1515] = n_Body_y[1515];
                c_Body_x[1516] = n_Body_x[1516];
                c_Body_y[1516] = n_Body_y[1516];
                c_Body_x[1517] = n_Body_x[1517];
                c_Body_y[1517] = n_Body_y[1517];
                c_Body_x[1518] = n_Body_x[1518];
                c_Body_y[1518] = n_Body_y[1518];
                c_Body_x[1519] = n_Body_x[1519];
                c_Body_y[1519] = n_Body_y[1519];
                c_Body_x[1520] = n_Body_x[1520];
                c_Body_y[1520] = n_Body_y[1520];
                c_Body_x[1521] = n_Body_x[1521];
                c_Body_y[1521] = n_Body_y[1521];
                c_Body_x[1522] = n_Body_x[1522];
                c_Body_y[1522] = n_Body_y[1522];
                c_Body_x[1523] = n_Body_x[1523];
                c_Body_y[1523] = n_Body_y[1523];
                c_Body_x[1524] = n_Body_x[1524];
                c_Body_y[1524] = n_Body_y[1524];
                c_Body_x[1525] = n_Body_x[1525];
                c_Body_y[1525] = n_Body_y[1525];
                c_Body_x[1526] = n_Body_x[1526];
                c_Body_y[1526] = n_Body_y[1526];
                c_Body_x[1527] = n_Body_x[1527];
                c_Body_y[1527] = n_Body_y[1527];
                c_Body_x[1528] = n_Body_x[1528];
                c_Body_y[1528] = n_Body_y[1528];
                c_Body_x[1529] = n_Body_x[1529];
                c_Body_y[1529] = n_Body_y[1529];
                c_Body_x[1530] = n_Body_x[1530];
                c_Body_y[1530] = n_Body_y[1530];
                c_Body_x[1531] = n_Body_x[1531];
                c_Body_y[1531] = n_Body_y[1531];
                c_Body_x[1532] = n_Body_x[1532];
                c_Body_y[1532] = n_Body_y[1532];
                c_Body_x[1533] = n_Body_x[1533];
                c_Body_y[1533] = n_Body_y[1533];
                c_Body_x[1534] = n_Body_x[1534];
                c_Body_y[1534] = n_Body_y[1534];
                c_Body_x[1535] = n_Body_x[1535];
                c_Body_y[1535] = n_Body_y[1535];
                c_Body_x[1536] = n_Body_x[1536];
                c_Body_y[1536] = n_Body_y[1536];
                c_Body_x[1537] = n_Body_x[1537];
                c_Body_y[1537] = n_Body_y[1537];
                c_Body_x[1538] = n_Body_x[1538];
                c_Body_y[1538] = n_Body_y[1538];
                c_Body_x[1539] = n_Body_x[1539];
                c_Body_y[1539] = n_Body_y[1539];
                c_Body_x[1540] = n_Body_x[1540];
                c_Body_y[1540] = n_Body_y[1540];
                c_Body_x[1541] = n_Body_x[1541];
                c_Body_y[1541] = n_Body_y[1541];
                c_Body_x[1542] = n_Body_x[1542];
                c_Body_y[1542] = n_Body_y[1542];
                c_Body_x[1543] = n_Body_x[1543];
                c_Body_y[1543] = n_Body_y[1543];
                c_Body_x[1544] = n_Body_x[1544];
                c_Body_y[1544] = n_Body_y[1544];
                c_Body_x[1545] = n_Body_x[1545];
                c_Body_y[1545] = n_Body_y[1545];
                c_Body_x[1546] = n_Body_x[1546];
                c_Body_y[1546] = n_Body_y[1546];
                c_Body_x[1547] = n_Body_x[1547];
                c_Body_y[1547] = n_Body_y[1547];
                c_Body_x[1548] = n_Body_x[1548];
                c_Body_y[1548] = n_Body_y[1548];
                c_Body_x[1549] = n_Body_x[1549];
                c_Body_y[1549] = n_Body_y[1549];
                c_Body_x[1550] = n_Body_x[1550];
                c_Body_y[1550] = n_Body_y[1550];
                c_Body_x[1551] = n_Body_x[1551];
                c_Body_y[1551] = n_Body_y[1551];
                c_Body_x[1552] = n_Body_x[1552];
                c_Body_y[1552] = n_Body_y[1552];
                c_Body_x[1553] = n_Body_x[1553];
                c_Body_y[1553] = n_Body_y[1553];
                c_Body_x[1554] = n_Body_x[1554];
                c_Body_y[1554] = n_Body_y[1554];
                c_Body_x[1555] = n_Body_x[1555];
                c_Body_y[1555] = n_Body_y[1555];
                c_Body_x[1556] = n_Body_x[1556];
                c_Body_y[1556] = n_Body_y[1556];
                c_Body_x[1557] = n_Body_x[1557];
                c_Body_y[1557] = n_Body_y[1557];
                c_Body_x[1558] = n_Body_x[1558];
                c_Body_y[1558] = n_Body_y[1558];
                c_Body_x[1559] = n_Body_x[1559];
                c_Body_y[1559] = n_Body_y[1559];
                c_Body_x[1560] = n_Body_x[1560];
                c_Body_y[1560] = n_Body_y[1560];
                c_Body_x[1561] = n_Body_x[1561];
                c_Body_y[1561] = n_Body_y[1561];
                c_Body_x[1562] = n_Body_x[1562];
                c_Body_y[1562] = n_Body_y[1562];
                c_Body_x[1563] = n_Body_x[1563];
                c_Body_y[1563] = n_Body_y[1563];
                c_Body_x[1564] = n_Body_x[1564];
                c_Body_y[1564] = n_Body_y[1564];
                c_Body_x[1565] = n_Body_x[1565];
                c_Body_y[1565] = n_Body_y[1565];
                c_Body_x[1566] = n_Body_x[1566];
                c_Body_y[1566] = n_Body_y[1566];
                c_Body_x[1567] = n_Body_x[1567];
                c_Body_y[1567] = n_Body_y[1567];
                c_Body_x[1568] = n_Body_x[1568];
                c_Body_y[1568] = n_Body_y[1568];
                c_Body_x[1569] = n_Body_x[1569];
                c_Body_y[1569] = n_Body_y[1569];
                c_Body_x[1570] = n_Body_x[1570];
                c_Body_y[1570] = n_Body_y[1570];
                c_Body_x[1571] = n_Body_x[1571];
                c_Body_y[1571] = n_Body_y[1571];
                c_Body_x[1572] = n_Body_x[1572];
                c_Body_y[1572] = n_Body_y[1572];
                c_Body_x[1573] = n_Body_x[1573];
                c_Body_y[1573] = n_Body_y[1573];
                c_Body_x[1574] = n_Body_x[1574];
                c_Body_y[1574] = n_Body_y[1574];
                c_Body_x[1575] = n_Body_x[1575];
                c_Body_y[1575] = n_Body_y[1575];
                c_Body_x[1576] = n_Body_x[1576];
                c_Body_y[1576] = n_Body_y[1576];
                c_Body_x[1577] = n_Body_x[1577];
                c_Body_y[1577] = n_Body_y[1577];
                c_Body_x[1578] = n_Body_x[1578];
                c_Body_y[1578] = n_Body_y[1578];
                c_Body_x[1579] = n_Body_x[1579];
                c_Body_y[1579] = n_Body_y[1579];
                c_Body_x[1580] = n_Body_x[1580];
                c_Body_y[1580] = n_Body_y[1580];
                c_Body_x[1581] = n_Body_x[1581];
                c_Body_y[1581] = n_Body_y[1581];
                c_Body_x[1582] = n_Body_x[1582];
                c_Body_y[1582] = n_Body_y[1582];
                c_Body_x[1583] = n_Body_x[1583];
                c_Body_y[1583] = n_Body_y[1583];
                c_Body_x[1584] = n_Body_x[1584];
                c_Body_y[1584] = n_Body_y[1584];
                c_Body_x[1585] = n_Body_x[1585];
                c_Body_y[1585] = n_Body_y[1585];
                c_Body_x[1586] = n_Body_x[1586];
                c_Body_y[1586] = n_Body_y[1586];
                c_Body_x[1587] = n_Body_x[1587];
                c_Body_y[1587] = n_Body_y[1587];
                c_Body_x[1588] = n_Body_x[1588];
                c_Body_y[1588] = n_Body_y[1588];
                c_Body_x[1589] = n_Body_x[1589];
                c_Body_y[1589] = n_Body_y[1589];
                c_Body_x[1590] = n_Body_x[1590];
                c_Body_y[1590] = n_Body_y[1590];
                c_Body_x[1591] = n_Body_x[1591];
                c_Body_y[1591] = n_Body_y[1591];
                c_Body_x[1592] = n_Body_x[1592];
                c_Body_y[1592] = n_Body_y[1592];
                c_Body_x[1593] = n_Body_x[1593];
                c_Body_y[1593] = n_Body_y[1593];
                c_Body_x[1594] = n_Body_x[1594];
                c_Body_y[1594] = n_Body_y[1594];
                c_Body_x[1595] = n_Body_x[1595];
                c_Body_y[1595] = n_Body_y[1595];
                c_Body_x[1596] = n_Body_x[1596];
                c_Body_y[1596] = n_Body_y[1596];
                c_Body_x[1597] = n_Body_x[1597];
                c_Body_y[1597] = n_Body_y[1597];
                c_Body_x[1598] = n_Body_x[1598];
                c_Body_y[1598] = n_Body_y[1598];
                c_Body_x[1599] = n_Body_x[1599];
                c_Body_y[1599] = n_Body_y[1599];
                c_Body_x[1600] = n_Body_x[1600];
                c_Body_y[1600] = n_Body_y[1600];
                c_Body_x[1601] = n_Body_x[1601];
                c_Body_y[1601] = n_Body_y[1601];
                c_Body_x[1602] = n_Body_x[1602];
                c_Body_y[1602] = n_Body_y[1602];
                c_Body_x[1603] = n_Body_x[1603];
                c_Body_y[1603] = n_Body_y[1603];
                c_Body_x[1604] = n_Body_x[1604];
                c_Body_y[1604] = n_Body_y[1604];
                c_Body_x[1605] = n_Body_x[1605];
                c_Body_y[1605] = n_Body_y[1605];
                c_Body_x[1606] = n_Body_x[1606];
                c_Body_y[1606] = n_Body_y[1606];
                c_Body_x[1607] = n_Body_x[1607];
                c_Body_y[1607] = n_Body_y[1607];
                c_Body_x[1608] = n_Body_x[1608];
                c_Body_y[1608] = n_Body_y[1608];
                c_Body_x[1609] = n_Body_x[1609];
                c_Body_y[1609] = n_Body_y[1609];
                c_Body_x[1610] = n_Body_x[1610];
                c_Body_y[1610] = n_Body_y[1610];
                c_Body_x[1611] = n_Body_x[1611];
                c_Body_y[1611] = n_Body_y[1611];
                c_Body_x[1612] = n_Body_x[1612];
                c_Body_y[1612] = n_Body_y[1612];
                c_Body_x[1613] = n_Body_x[1613];
                c_Body_y[1613] = n_Body_y[1613];
                c_Body_x[1614] = n_Body_x[1614];
                c_Body_y[1614] = n_Body_y[1614];
                c_Body_x[1615] = n_Body_x[1615];
                c_Body_y[1615] = n_Body_y[1615];
                c_Body_x[1616] = n_Body_x[1616];
                c_Body_y[1616] = n_Body_y[1616];
                c_Body_x[1617] = n_Body_x[1617];
                c_Body_y[1617] = n_Body_y[1617];
                c_Body_x[1618] = n_Body_x[1618];
                c_Body_y[1618] = n_Body_y[1618];
                c_Body_x[1619] = n_Body_x[1619];
                c_Body_y[1619] = n_Body_y[1619];
                c_Body_x[1620] = n_Body_x[1620];
                c_Body_y[1620] = n_Body_y[1620];
                c_Body_x[1621] = n_Body_x[1621];
                c_Body_y[1621] = n_Body_y[1621];
                c_Body_x[1622] = n_Body_x[1622];
                c_Body_y[1622] = n_Body_y[1622];
                c_Body_x[1623] = n_Body_x[1623];
                c_Body_y[1623] = n_Body_y[1623];
                c_Body_x[1624] = n_Body_x[1624];
                c_Body_y[1624] = n_Body_y[1624];
                c_Body_x[1625] = n_Body_x[1625];
                c_Body_y[1625] = n_Body_y[1625];
                c_Body_x[1626] = n_Body_x[1626];
                c_Body_y[1626] = n_Body_y[1626];
                c_Body_x[1627] = n_Body_x[1627];
                c_Body_y[1627] = n_Body_y[1627];
                c_Body_x[1628] = n_Body_x[1628];
                c_Body_y[1628] = n_Body_y[1628];
                c_Body_x[1629] = n_Body_x[1629];
                c_Body_y[1629] = n_Body_y[1629];
                c_Body_x[1630] = n_Body_x[1630];
                c_Body_y[1630] = n_Body_y[1630];
                c_Body_x[1631] = n_Body_x[1631];
                c_Body_y[1631] = n_Body_y[1631];
                c_Body_x[1632] = n_Body_x[1632];
                c_Body_y[1632] = n_Body_y[1632];
                c_Body_x[1633] = n_Body_x[1633];
                c_Body_y[1633] = n_Body_y[1633];
                c_Body_x[1634] = n_Body_x[1634];
                c_Body_y[1634] = n_Body_y[1634];
                c_Body_x[1635] = n_Body_x[1635];
                c_Body_y[1635] = n_Body_y[1635];
                c_Body_x[1636] = n_Body_x[1636];
                c_Body_y[1636] = n_Body_y[1636];
                c_Body_x[1637] = n_Body_x[1637];
                c_Body_y[1637] = n_Body_y[1637];
                c_Body_x[1638] = n_Body_x[1638];
                c_Body_y[1638] = n_Body_y[1638];
                c_Body_x[1639] = n_Body_x[1639];
                c_Body_y[1639] = n_Body_y[1639];
                c_Body_x[1640] = n_Body_x[1640];
                c_Body_y[1640] = n_Body_y[1640];
                c_Body_x[1641] = n_Body_x[1641];
                c_Body_y[1641] = n_Body_y[1641];
                c_Body_x[1642] = n_Body_x[1642];
                c_Body_y[1642] = n_Body_y[1642];
                c_Body_x[1643] = n_Body_x[1643];
                c_Body_y[1643] = n_Body_y[1643];
                c_Body_x[1644] = n_Body_x[1644];
                c_Body_y[1644] = n_Body_y[1644];
                c_Body_x[1645] = n_Body_x[1645];
                c_Body_y[1645] = n_Body_y[1645];
                c_Body_x[1646] = n_Body_x[1646];
                c_Body_y[1646] = n_Body_y[1646];
                c_Body_x[1647] = n_Body_x[1647];
                c_Body_y[1647] = n_Body_y[1647];
                c_Body_x[1648] = n_Body_x[1648];
                c_Body_y[1648] = n_Body_y[1648];
                c_Body_x[1649] = n_Body_x[1649];
                c_Body_y[1649] = n_Body_y[1649];
                c_Body_x[1650] = n_Body_x[1650];
                c_Body_y[1650] = n_Body_y[1650];
                c_Body_x[1651] = n_Body_x[1651];
                c_Body_y[1651] = n_Body_y[1651];
                c_Body_x[1652] = n_Body_x[1652];
                c_Body_y[1652] = n_Body_y[1652];
                c_Body_x[1653] = n_Body_x[1653];
                c_Body_y[1653] = n_Body_y[1653];
                c_Body_x[1654] = n_Body_x[1654];
                c_Body_y[1654] = n_Body_y[1654];
                c_Body_x[1655] = n_Body_x[1655];
                c_Body_y[1655] = n_Body_y[1655];
                c_Body_x[1656] = n_Body_x[1656];
                c_Body_y[1656] = n_Body_y[1656];
                c_Body_x[1657] = n_Body_x[1657];
                c_Body_y[1657] = n_Body_y[1657];
                c_Body_x[1658] = n_Body_x[1658];
                c_Body_y[1658] = n_Body_y[1658];
                c_Body_x[1659] = n_Body_x[1659];
                c_Body_y[1659] = n_Body_y[1659];
                c_Body_x[1660] = n_Body_x[1660];
                c_Body_y[1660] = n_Body_y[1660];
                c_Body_x[1661] = n_Body_x[1661];
                c_Body_y[1661] = n_Body_y[1661];
                c_Body_x[1662] = n_Body_x[1662];
                c_Body_y[1662] = n_Body_y[1662];
                c_Body_x[1663] = n_Body_x[1663];
                c_Body_y[1663] = n_Body_y[1663];
                c_Body_x[1664] = n_Body_x[1664];
                c_Body_y[1664] = n_Body_y[1664];
                c_Body_x[1665] = n_Body_x[1665];
                c_Body_y[1665] = n_Body_y[1665];
                c_Body_x[1666] = n_Body_x[1666];
                c_Body_y[1666] = n_Body_y[1666];
                c_Body_x[1667] = n_Body_x[1667];
                c_Body_y[1667] = n_Body_y[1667];
                c_Body_x[1668] = n_Body_x[1668];
                c_Body_y[1668] = n_Body_y[1668];
                c_Body_x[1669] = n_Body_x[1669];
                c_Body_y[1669] = n_Body_y[1669];
                c_Body_x[1670] = n_Body_x[1670];
                c_Body_y[1670] = n_Body_y[1670];
                c_Body_x[1671] = n_Body_x[1671];
                c_Body_y[1671] = n_Body_y[1671];
                c_Body_x[1672] = n_Body_x[1672];
                c_Body_y[1672] = n_Body_y[1672];
                c_Body_x[1673] = n_Body_x[1673];
                c_Body_y[1673] = n_Body_y[1673];
                c_Body_x[1674] = n_Body_x[1674];
                c_Body_y[1674] = n_Body_y[1674];
                c_Body_x[1675] = n_Body_x[1675];
                c_Body_y[1675] = n_Body_y[1675];
                c_Body_x[1676] = n_Body_x[1676];
                c_Body_y[1676] = n_Body_y[1676];
                c_Body_x[1677] = n_Body_x[1677];
                c_Body_y[1677] = n_Body_y[1677];
                c_Body_x[1678] = n_Body_x[1678];
                c_Body_y[1678] = n_Body_y[1678];
                c_Body_x[1679] = n_Body_x[1679];
                c_Body_y[1679] = n_Body_y[1679];
                c_Body_x[1680] = n_Body_x[1680];
                c_Body_y[1680] = n_Body_y[1680];
                c_Body_x[1681] = n_Body_x[1681];
                c_Body_y[1681] = n_Body_y[1681];
                c_Body_x[1682] = n_Body_x[1682];
                c_Body_y[1682] = n_Body_y[1682];
                c_Body_x[1683] = n_Body_x[1683];
                c_Body_y[1683] = n_Body_y[1683];
                c_Body_x[1684] = n_Body_x[1684];
                c_Body_y[1684] = n_Body_y[1684];
                c_Body_x[1685] = n_Body_x[1685];
                c_Body_y[1685] = n_Body_y[1685];
                c_Body_x[1686] = n_Body_x[1686];
                c_Body_y[1686] = n_Body_y[1686];
                c_Body_x[1687] = n_Body_x[1687];
                c_Body_y[1687] = n_Body_y[1687];
                c_Body_x[1688] = n_Body_x[1688];
                c_Body_y[1688] = n_Body_y[1688];
                c_Body_x[1689] = n_Body_x[1689];
                c_Body_y[1689] = n_Body_y[1689];
                c_Body_x[1690] = n_Body_x[1690];
                c_Body_y[1690] = n_Body_y[1690];
                c_Body_x[1691] = n_Body_x[1691];
                c_Body_y[1691] = n_Body_y[1691];
                c_Body_x[1692] = n_Body_x[1692];
                c_Body_y[1692] = n_Body_y[1692];
                c_Body_x[1693] = n_Body_x[1693];
                c_Body_y[1693] = n_Body_y[1693];
                c_Body_x[1694] = n_Body_x[1694];
                c_Body_y[1694] = n_Body_y[1694];
                c_Body_x[1695] = n_Body_x[1695];
                c_Body_y[1695] = n_Body_y[1695];
                c_Body_x[1696] = n_Body_x[1696];
                c_Body_y[1696] = n_Body_y[1696];
                c_Body_x[1697] = n_Body_x[1697];
                c_Body_y[1697] = n_Body_y[1697];
                c_Body_x[1698] = n_Body_x[1698];
                c_Body_y[1698] = n_Body_y[1698];
                c_Body_x[1699] = n_Body_x[1699];
                c_Body_y[1699] = n_Body_y[1699];
                c_Body_x[1700] = n_Body_x[1700];
                c_Body_y[1700] = n_Body_y[1700];
                c_Body_x[1701] = n_Body_x[1701];
                c_Body_y[1701] = n_Body_y[1701];
                c_Body_x[1702] = n_Body_x[1702];
                c_Body_y[1702] = n_Body_y[1702];
                c_Body_x[1703] = n_Body_x[1703];
                c_Body_y[1703] = n_Body_y[1703];
                c_Body_x[1704] = n_Body_x[1704];
                c_Body_y[1704] = n_Body_y[1704];
                c_Body_x[1705] = n_Body_x[1705];
                c_Body_y[1705] = n_Body_y[1705];
                c_Body_x[1706] = n_Body_x[1706];
                c_Body_y[1706] = n_Body_y[1706];
                c_Body_x[1707] = n_Body_x[1707];
                c_Body_y[1707] = n_Body_y[1707];
                c_Body_x[1708] = n_Body_x[1708];
                c_Body_y[1708] = n_Body_y[1708];
                c_Body_x[1709] = n_Body_x[1709];
                c_Body_y[1709] = n_Body_y[1709];
                c_Body_x[1710] = n_Body_x[1710];
                c_Body_y[1710] = n_Body_y[1710];
                c_Body_x[1711] = n_Body_x[1711];
                c_Body_y[1711] = n_Body_y[1711];
                c_Body_x[1712] = n_Body_x[1712];
                c_Body_y[1712] = n_Body_y[1712];
                c_Body_x[1713] = n_Body_x[1713];
                c_Body_y[1713] = n_Body_y[1713];
                c_Body_x[1714] = n_Body_x[1714];
                c_Body_y[1714] = n_Body_y[1714];
                c_Body_x[1715] = n_Body_x[1715];
                c_Body_y[1715] = n_Body_y[1715];
                c_Body_x[1716] = n_Body_x[1716];
                c_Body_y[1716] = n_Body_y[1716];
                c_Body_x[1717] = n_Body_x[1717];
                c_Body_y[1717] = n_Body_y[1717];
                c_Body_x[1718] = n_Body_x[1718];
                c_Body_y[1718] = n_Body_y[1718];
                c_Body_x[1719] = n_Body_x[1719];
                c_Body_y[1719] = n_Body_y[1719];
                c_Body_x[1720] = n_Body_x[1720];
                c_Body_y[1720] = n_Body_y[1720];
                c_Body_x[1721] = n_Body_x[1721];
                c_Body_y[1721] = n_Body_y[1721];
                c_Body_x[1722] = n_Body_x[1722];
                c_Body_y[1722] = n_Body_y[1722];
                c_Body_x[1723] = n_Body_x[1723];
                c_Body_y[1723] = n_Body_y[1723];
                c_Body_x[1724] = n_Body_x[1724];
                c_Body_y[1724] = n_Body_y[1724];
                c_Body_x[1725] = n_Body_x[1725];
                c_Body_y[1725] = n_Body_y[1725];
                c_Body_x[1726] = n_Body_x[1726];
                c_Body_y[1726] = n_Body_y[1726];
                c_Body_x[1727] = n_Body_x[1727];
                c_Body_y[1727] = n_Body_y[1727];
                c_Body_x[1728] = n_Body_x[1728];
                c_Body_y[1728] = n_Body_y[1728];
                c_Body_x[1729] = n_Body_x[1729];
                c_Body_y[1729] = n_Body_y[1729];
                c_Body_x[1730] = n_Body_x[1730];
                c_Body_y[1730] = n_Body_y[1730];
                c_Body_x[1731] = n_Body_x[1731];
                c_Body_y[1731] = n_Body_y[1731];
                c_Body_x[1732] = n_Body_x[1732];
                c_Body_y[1732] = n_Body_y[1732];
                c_Body_x[1733] = n_Body_x[1733];
                c_Body_y[1733] = n_Body_y[1733];
                c_Body_x[1734] = n_Body_x[1734];
                c_Body_y[1734] = n_Body_y[1734];
                c_Body_x[1735] = n_Body_x[1735];
                c_Body_y[1735] = n_Body_y[1735];
                c_Body_x[1736] = n_Body_x[1736];
                c_Body_y[1736] = n_Body_y[1736];
                c_Body_x[1737] = n_Body_x[1737];
                c_Body_y[1737] = n_Body_y[1737];
                c_Body_x[1738] = n_Body_x[1738];
                c_Body_y[1738] = n_Body_y[1738];
                c_Body_x[1739] = n_Body_x[1739];
                c_Body_y[1739] = n_Body_y[1739];
                c_Body_x[1740] = n_Body_x[1740];
                c_Body_y[1740] = n_Body_y[1740];
                c_Body_x[1741] = n_Body_x[1741];
                c_Body_y[1741] = n_Body_y[1741];
                c_Body_x[1742] = n_Body_x[1742];
                c_Body_y[1742] = n_Body_y[1742];
                c_Body_x[1743] = n_Body_x[1743];
                c_Body_y[1743] = n_Body_y[1743];
                c_Body_x[1744] = n_Body_x[1744];
                c_Body_y[1744] = n_Body_y[1744];
                c_Body_x[1745] = n_Body_x[1745];
                c_Body_y[1745] = n_Body_y[1745];
                c_Body_x[1746] = n_Body_x[1746];
                c_Body_y[1746] = n_Body_y[1746];
                c_Body_x[1747] = n_Body_x[1747];
                c_Body_y[1747] = n_Body_y[1747];
                c_Body_x[1748] = n_Body_x[1748];
                c_Body_y[1748] = n_Body_y[1748];
                c_Body_x[1749] = n_Body_x[1749];
                c_Body_y[1749] = n_Body_y[1749];
                c_Body_x[1750] = n_Body_x[1750];
                c_Body_y[1750] = n_Body_y[1750];
                c_Body_x[1751] = n_Body_x[1751];
                c_Body_y[1751] = n_Body_y[1751];
                c_Body_x[1752] = n_Body_x[1752];
                c_Body_y[1752] = n_Body_y[1752];
                c_Body_x[1753] = n_Body_x[1753];
                c_Body_y[1753] = n_Body_y[1753];
                c_Body_x[1754] = n_Body_x[1754];
                c_Body_y[1754] = n_Body_y[1754];
                c_Body_x[1755] = n_Body_x[1755];
                c_Body_y[1755] = n_Body_y[1755];
                c_Body_x[1756] = n_Body_x[1756];
                c_Body_y[1756] = n_Body_y[1756];
                c_Body_x[1757] = n_Body_x[1757];
                c_Body_y[1757] = n_Body_y[1757];
                c_Body_x[1758] = n_Body_x[1758];
                c_Body_y[1758] = n_Body_y[1758];
                c_Body_x[1759] = n_Body_x[1759];
                c_Body_y[1759] = n_Body_y[1759];
                c_Body_x[1760] = n_Body_x[1760];
                c_Body_y[1760] = n_Body_y[1760];
                c_Body_x[1761] = n_Body_x[1761];
                c_Body_y[1761] = n_Body_y[1761];
                c_Body_x[1762] = n_Body_x[1762];
                c_Body_y[1762] = n_Body_y[1762];
                c_Body_x[1763] = n_Body_x[1763];
                c_Body_y[1763] = n_Body_y[1763];
                c_Body_x[1764] = n_Body_x[1764];
                c_Body_y[1764] = n_Body_y[1764];
                c_Body_x[1765] = n_Body_x[1765];
                c_Body_y[1765] = n_Body_y[1765];
                c_Body_x[1766] = n_Body_x[1766];
                c_Body_y[1766] = n_Body_y[1766];
                c_Body_x[1767] = n_Body_x[1767];
                c_Body_y[1767] = n_Body_y[1767];
                c_Body_x[1768] = n_Body_x[1768];
                c_Body_y[1768] = n_Body_y[1768];
                c_Body_x[1769] = n_Body_x[1769];
                c_Body_y[1769] = n_Body_y[1769];
                c_Body_x[1770] = n_Body_x[1770];
                c_Body_y[1770] = n_Body_y[1770];
                c_Body_x[1771] = n_Body_x[1771];
                c_Body_y[1771] = n_Body_y[1771];
                c_Body_x[1772] = n_Body_x[1772];
                c_Body_y[1772] = n_Body_y[1772];
                c_Body_x[1773] = n_Body_x[1773];
                c_Body_y[1773] = n_Body_y[1773];
                c_Body_x[1774] = n_Body_x[1774];
                c_Body_y[1774] = n_Body_y[1774];
                c_Body_x[1775] = n_Body_x[1775];
                c_Body_y[1775] = n_Body_y[1775];
                c_Body_x[1776] = n_Body_x[1776];
                c_Body_y[1776] = n_Body_y[1776];
                c_Body_x[1777] = n_Body_x[1777];
                c_Body_y[1777] = n_Body_y[1777];
                c_Body_x[1778] = n_Body_x[1778];
                c_Body_y[1778] = n_Body_y[1778];
                c_Body_x[1779] = n_Body_x[1779];
                c_Body_y[1779] = n_Body_y[1779];
                c_Body_x[1780] = n_Body_x[1780];
                c_Body_y[1780] = n_Body_y[1780];
                c_Body_x[1781] = n_Body_x[1781];
                c_Body_y[1781] = n_Body_y[1781];
                c_Body_x[1782] = n_Body_x[1782];
                c_Body_y[1782] = n_Body_y[1782];
                c_Body_x[1783] = n_Body_x[1783];
                c_Body_y[1783] = n_Body_y[1783];
                c_Body_x[1784] = n_Body_x[1784];
                c_Body_y[1784] = n_Body_y[1784];
                c_Body_x[1785] = n_Body_x[1785];
                c_Body_y[1785] = n_Body_y[1785];
                c_Body_x[1786] = n_Body_x[1786];
                c_Body_y[1786] = n_Body_y[1786];
                c_Body_x[1787] = n_Body_x[1787];
                c_Body_y[1787] = n_Body_y[1787];
                c_Body_x[1788] = n_Body_x[1788];
                c_Body_y[1788] = n_Body_y[1788];
                c_Body_x[1789] = n_Body_x[1789];
                c_Body_y[1789] = n_Body_y[1789];
                c_Body_x[1790] = n_Body_x[1790];
                c_Body_y[1790] = n_Body_y[1790];
                c_Body_x[1791] = n_Body_x[1791];
                c_Body_y[1791] = n_Body_y[1791];
                c_Body_x[1792] = n_Body_x[1792];
                c_Body_y[1792] = n_Body_y[1792];
                c_Body_x[1793] = n_Body_x[1793];
                c_Body_y[1793] = n_Body_y[1793];
                c_Body_x[1794] = n_Body_x[1794];
                c_Body_y[1794] = n_Body_y[1794];
                c_Body_x[1795] = n_Body_x[1795];
                c_Body_y[1795] = n_Body_y[1795];
                c_Body_x[1796] = n_Body_x[1796];
                c_Body_y[1796] = n_Body_y[1796];
                c_Body_x[1797] = n_Body_x[1797];
                c_Body_y[1797] = n_Body_y[1797];
                c_Body_x[1798] = n_Body_x[1798];
                c_Body_y[1798] = n_Body_y[1798];
                c_Body_x[1799] = n_Body_x[1799];
                c_Body_y[1799] = n_Body_y[1799];
                c_Body_x[1800] = n_Body_x[1800];
                c_Body_y[1800] = n_Body_y[1800];
                c_Body_x[1801] = n_Body_x[1801];
                c_Body_y[1801] = n_Body_y[1801];
                c_Body_x[1802] = n_Body_x[1802];
                c_Body_y[1802] = n_Body_y[1802];
                c_Body_x[1803] = n_Body_x[1803];
                c_Body_y[1803] = n_Body_y[1803];
                c_Body_x[1804] = n_Body_x[1804];
                c_Body_y[1804] = n_Body_y[1804];
                c_Body_x[1805] = n_Body_x[1805];
                c_Body_y[1805] = n_Body_y[1805];
                c_Body_x[1806] = n_Body_x[1806];
                c_Body_y[1806] = n_Body_y[1806];
                c_Body_x[1807] = n_Body_x[1807];
                c_Body_y[1807] = n_Body_y[1807];
                c_Body_x[1808] = n_Body_x[1808];
                c_Body_y[1808] = n_Body_y[1808];
                c_Body_x[1809] = n_Body_x[1809];
                c_Body_y[1809] = n_Body_y[1809];
                c_Body_x[1810] = n_Body_x[1810];
                c_Body_y[1810] = n_Body_y[1810];
                c_Body_x[1811] = n_Body_x[1811];
                c_Body_y[1811] = n_Body_y[1811];
                c_Body_x[1812] = n_Body_x[1812];
                c_Body_y[1812] = n_Body_y[1812];
                c_Body_x[1813] = n_Body_x[1813];
                c_Body_y[1813] = n_Body_y[1813];
                c_Body_x[1814] = n_Body_x[1814];
                c_Body_y[1814] = n_Body_y[1814];
                c_Body_x[1815] = n_Body_x[1815];
                c_Body_y[1815] = n_Body_y[1815];
                c_Body_x[1816] = n_Body_x[1816];
                c_Body_y[1816] = n_Body_y[1816];
                c_Body_x[1817] = n_Body_x[1817];
                c_Body_y[1817] = n_Body_y[1817];
                c_Body_x[1818] = n_Body_x[1818];
                c_Body_y[1818] = n_Body_y[1818];
                c_Body_x[1819] = n_Body_x[1819];
                c_Body_y[1819] = n_Body_y[1819];
                c_Body_x[1820] = n_Body_x[1820];
                c_Body_y[1820] = n_Body_y[1820];
                c_Body_x[1821] = n_Body_x[1821];
                c_Body_y[1821] = n_Body_y[1821];
                c_Body_x[1822] = n_Body_x[1822];
                c_Body_y[1822] = n_Body_y[1822];
                c_Body_x[1823] = n_Body_x[1823];
                c_Body_y[1823] = n_Body_y[1823];
                c_Body_x[1824] = n_Body_x[1824];
                c_Body_y[1824] = n_Body_y[1824];
                c_Body_x[1825] = n_Body_x[1825];
                c_Body_y[1825] = n_Body_y[1825];
                c_Body_x[1826] = n_Body_x[1826];
                c_Body_y[1826] = n_Body_y[1826];
                c_Body_x[1827] = n_Body_x[1827];
                c_Body_y[1827] = n_Body_y[1827];
                c_Body_x[1828] = n_Body_x[1828];
                c_Body_y[1828] = n_Body_y[1828];
                c_Body_x[1829] = n_Body_x[1829];
                c_Body_y[1829] = n_Body_y[1829];
                c_Body_x[1830] = n_Body_x[1830];
                c_Body_y[1830] = n_Body_y[1830];
                c_Body_x[1831] = n_Body_x[1831];
                c_Body_y[1831] = n_Body_y[1831];
                c_Body_x[1832] = n_Body_x[1832];
                c_Body_y[1832] = n_Body_y[1832];
                c_Body_x[1833] = n_Body_x[1833];
                c_Body_y[1833] = n_Body_y[1833];
                c_Body_x[1834] = n_Body_x[1834];
                c_Body_y[1834] = n_Body_y[1834];
                c_Body_x[1835] = n_Body_x[1835];
                c_Body_y[1835] = n_Body_y[1835];
                c_Body_x[1836] = n_Body_x[1836];
                c_Body_y[1836] = n_Body_y[1836];
                c_Body_x[1837] = n_Body_x[1837];
                c_Body_y[1837] = n_Body_y[1837];
                c_Body_x[1838] = n_Body_x[1838];
                c_Body_y[1838] = n_Body_y[1838];
                c_Body_x[1839] = n_Body_x[1839];
                c_Body_y[1839] = n_Body_y[1839];
                c_Body_x[1840] = n_Body_x[1840];
                c_Body_y[1840] = n_Body_y[1840];
                c_Body_x[1841] = n_Body_x[1841];
                c_Body_y[1841] = n_Body_y[1841];
                c_Body_x[1842] = n_Body_x[1842];
                c_Body_y[1842] = n_Body_y[1842];
                c_Body_x[1843] = n_Body_x[1843];
                c_Body_y[1843] = n_Body_y[1843];
                c_Body_x[1844] = n_Body_x[1844];
                c_Body_y[1844] = n_Body_y[1844];
                c_Body_x[1845] = n_Body_x[1845];
                c_Body_y[1845] = n_Body_y[1845];
                c_Body_x[1846] = n_Body_x[1846];
                c_Body_y[1846] = n_Body_y[1846];
                c_Body_x[1847] = n_Body_x[1847];
                c_Body_y[1847] = n_Body_y[1847];
                c_Body_x[1848] = n_Body_x[1848];
                c_Body_y[1848] = n_Body_y[1848];
                c_Body_x[1849] = n_Body_x[1849];
                c_Body_y[1849] = n_Body_y[1849];
                c_Body_x[1850] = n_Body_x[1850];
                c_Body_y[1850] = n_Body_y[1850];
                c_Body_x[1851] = n_Body_x[1851];
                c_Body_y[1851] = n_Body_y[1851];
                c_Body_x[1852] = n_Body_x[1852];
                c_Body_y[1852] = n_Body_y[1852];
                c_Body_x[1853] = n_Body_x[1853];
                c_Body_y[1853] = n_Body_y[1853];
                c_Body_x[1854] = n_Body_x[1854];
                c_Body_y[1854] = n_Body_y[1854];
                c_Body_x[1855] = n_Body_x[1855];
                c_Body_y[1855] = n_Body_y[1855];
                c_Body_x[1856] = n_Body_x[1856];
                c_Body_y[1856] = n_Body_y[1856];
                c_Body_x[1857] = n_Body_x[1857];
                c_Body_y[1857] = n_Body_y[1857];
                c_Body_x[1858] = n_Body_x[1858];
                c_Body_y[1858] = n_Body_y[1858];
                c_Body_x[1859] = n_Body_x[1859];
                c_Body_y[1859] = n_Body_y[1859];
                c_Body_x[1860] = n_Body_x[1860];
                c_Body_y[1860] = n_Body_y[1860];
                c_Body_x[1861] = n_Body_x[1861];
                c_Body_y[1861] = n_Body_y[1861];
                c_Body_x[1862] = n_Body_x[1862];
                c_Body_y[1862] = n_Body_y[1862];
                c_Body_x[1863] = n_Body_x[1863];
                c_Body_y[1863] = n_Body_y[1863];
                c_Body_x[1864] = n_Body_x[1864];
                c_Body_y[1864] = n_Body_y[1864];
                c_Body_x[1865] = n_Body_x[1865];
                c_Body_y[1865] = n_Body_y[1865];
                c_Body_x[1866] = n_Body_x[1866];
                c_Body_y[1866] = n_Body_y[1866];
                c_Body_x[1867] = n_Body_x[1867];
                c_Body_y[1867] = n_Body_y[1867];
                c_Body_x[1868] = n_Body_x[1868];
                c_Body_y[1868] = n_Body_y[1868];
                c_Body_x[1869] = n_Body_x[1869];
                c_Body_y[1869] = n_Body_y[1869];
                c_Body_x[1870] = n_Body_x[1870];
                c_Body_y[1870] = n_Body_y[1870];
                c_Body_x[1871] = n_Body_x[1871];
                c_Body_y[1871] = n_Body_y[1871];
                c_Body_x[1872] = n_Body_x[1872];
                c_Body_y[1872] = n_Body_y[1872];
                c_Body_x[1873] = n_Body_x[1873];
                c_Body_y[1873] = n_Body_y[1873];
                c_Body_x[1874] = n_Body_x[1874];
                c_Body_y[1874] = n_Body_y[1874];
                c_Body_x[1875] = n_Body_x[1875];
                c_Body_y[1875] = n_Body_y[1875];
                c_Body_x[1876] = n_Body_x[1876];
                c_Body_y[1876] = n_Body_y[1876];
                c_Body_x[1877] = n_Body_x[1877];
                c_Body_y[1877] = n_Body_y[1877];
                c_Body_x[1878] = n_Body_x[1878];
                c_Body_y[1878] = n_Body_y[1878];
                c_Body_x[1879] = n_Body_x[1879];
                c_Body_y[1879] = n_Body_y[1879];
                c_Body_x[1880] = n_Body_x[1880];
                c_Body_y[1880] = n_Body_y[1880];
                c_Body_x[1881] = n_Body_x[1881];
                c_Body_y[1881] = n_Body_y[1881];
                c_Body_x[1882] = n_Body_x[1882];
                c_Body_y[1882] = n_Body_y[1882];
                c_Body_x[1883] = n_Body_x[1883];
                c_Body_y[1883] = n_Body_y[1883];
                c_Body_x[1884] = n_Body_x[1884];
                c_Body_y[1884] = n_Body_y[1884];
                c_Body_x[1885] = n_Body_x[1885];
                c_Body_y[1885] = n_Body_y[1885];
                c_Body_x[1886] = n_Body_x[1886];
                c_Body_y[1886] = n_Body_y[1886];
                c_Body_x[1887] = n_Body_x[1887];
                c_Body_y[1887] = n_Body_y[1887];
                c_Body_x[1888] = n_Body_x[1888];
                c_Body_y[1888] = n_Body_y[1888];
                c_Body_x[1889] = n_Body_x[1889];
                c_Body_y[1889] = n_Body_y[1889];
                c_Body_x[1890] = n_Body_x[1890];
                c_Body_y[1890] = n_Body_y[1890];
                c_Body_x[1891] = n_Body_x[1891];
                c_Body_y[1891] = n_Body_y[1891];
                c_Body_x[1892] = n_Body_x[1892];
                c_Body_y[1892] = n_Body_y[1892];
                c_Body_x[1893] = n_Body_x[1893];
                c_Body_y[1893] = n_Body_y[1893];
                c_Body_x[1894] = n_Body_x[1894];
                c_Body_y[1894] = n_Body_y[1894];
                c_Body_x[1895] = n_Body_x[1895];
                c_Body_y[1895] = n_Body_y[1895];
                c_Body_x[1896] = n_Body_x[1896];
                c_Body_y[1896] = n_Body_y[1896];
                c_Body_x[1897] = n_Body_x[1897];
                c_Body_y[1897] = n_Body_y[1897];
                c_Body_x[1898] = n_Body_x[1898];
                c_Body_y[1898] = n_Body_y[1898];
                c_Body_x[1899] = n_Body_x[1899];
                c_Body_y[1899] = n_Body_y[1899];
                c_Body_x[1900] = n_Body_x[1900];
                c_Body_y[1900] = n_Body_y[1900];
                c_Body_x[1901] = n_Body_x[1901];
                c_Body_y[1901] = n_Body_y[1901];
                c_Body_x[1902] = n_Body_x[1902];
                c_Body_y[1902] = n_Body_y[1902];
                c_Body_x[1903] = n_Body_x[1903];
                c_Body_y[1903] = n_Body_y[1903];
                c_Body_x[1904] = n_Body_x[1904];
                c_Body_y[1904] = n_Body_y[1904];
                c_Body_x[1905] = n_Body_x[1905];
                c_Body_y[1905] = n_Body_y[1905];
                c_Body_x[1906] = n_Body_x[1906];
                c_Body_y[1906] = n_Body_y[1906];
                c_Body_x[1907] = n_Body_x[1907];
                c_Body_y[1907] = n_Body_y[1907];
                c_Body_x[1908] = n_Body_x[1908];
                c_Body_y[1908] = n_Body_y[1908];
                c_Body_x[1909] = n_Body_x[1909];
                c_Body_y[1909] = n_Body_y[1909];
                c_Body_x[1910] = n_Body_x[1910];
                c_Body_y[1910] = n_Body_y[1910];
                c_Body_x[1911] = n_Body_x[1911];
                c_Body_y[1911] = n_Body_y[1911];
                c_Body_x[1912] = n_Body_x[1912];
                c_Body_y[1912] = n_Body_y[1912];
                c_Body_x[1913] = n_Body_x[1913];
                c_Body_y[1913] = n_Body_y[1913];
                c_Body_x[1914] = n_Body_x[1914];
                c_Body_y[1914] = n_Body_y[1914];
                c_Body_x[1915] = n_Body_x[1915];
                c_Body_y[1915] = n_Body_y[1915];
                c_Body_x[1916] = n_Body_x[1916];
                c_Body_y[1916] = n_Body_y[1916];
                c_Body_x[1917] = n_Body_x[1917];
                c_Body_y[1917] = n_Body_y[1917];
                c_Body_x[1918] = n_Body_x[1918];
                c_Body_y[1918] = n_Body_y[1918];
                c_Body_x[1919] = n_Body_x[1919];
                c_Body_y[1919] = n_Body_y[1919];
                c_Body_x[1920] = n_Body_x[1920];
                c_Body_y[1920] = n_Body_y[1920];
                c_Body_x[1921] = n_Body_x[1921];
                c_Body_y[1921] = n_Body_y[1921];
                c_Body_x[1922] = n_Body_x[1922];
                c_Body_y[1922] = n_Body_y[1922];
                c_Body_x[1923] = n_Body_x[1923];
                c_Body_y[1923] = n_Body_y[1923];
                c_Body_x[1924] = n_Body_x[1924];
                c_Body_y[1924] = n_Body_y[1924];
                c_Body_x[1925] = n_Body_x[1925];
                c_Body_y[1925] = n_Body_y[1925];
                c_Body_x[1926] = n_Body_x[1926];
                c_Body_y[1926] = n_Body_y[1926];
                c_Body_x[1927] = n_Body_x[1927];
                c_Body_y[1927] = n_Body_y[1927];
                c_Body_x[1928] = n_Body_x[1928];
                c_Body_y[1928] = n_Body_y[1928];
                c_Body_x[1929] = n_Body_x[1929];
                c_Body_y[1929] = n_Body_y[1929];
                c_Body_x[1930] = n_Body_x[1930];
                c_Body_y[1930] = n_Body_y[1930];
                c_Body_x[1931] = n_Body_x[1931];
                c_Body_y[1931] = n_Body_y[1931];
                c_Body_x[1932] = n_Body_x[1932];
                c_Body_y[1932] = n_Body_y[1932];
                c_Body_x[1933] = n_Body_x[1933];
                c_Body_y[1933] = n_Body_y[1933];
                c_Body_x[1934] = n_Body_x[1934];
                c_Body_y[1934] = n_Body_y[1934];
                c_Body_x[1935] = n_Body_x[1935];
                c_Body_y[1935] = n_Body_y[1935];
                c_Body_x[1936] = n_Body_x[1936];
                c_Body_y[1936] = n_Body_y[1936];
                c_Body_x[1937] = n_Body_x[1937];
                c_Body_y[1937] = n_Body_y[1937];
                c_Body_x[1938] = n_Body_x[1938];
                c_Body_y[1938] = n_Body_y[1938];
                c_Body_x[1939] = n_Body_x[1939];
                c_Body_y[1939] = n_Body_y[1939];
                c_Body_x[1940] = n_Body_x[1940];
                c_Body_y[1940] = n_Body_y[1940];
                c_Body_x[1941] = n_Body_x[1941];
                c_Body_y[1941] = n_Body_y[1941];
                c_Body_x[1942] = n_Body_x[1942];
                c_Body_y[1942] = n_Body_y[1942];
                c_Body_x[1943] = n_Body_x[1943];
                c_Body_y[1943] = n_Body_y[1943];
                c_Body_x[1944] = n_Body_x[1944];
                c_Body_y[1944] = n_Body_y[1944];
                c_Body_x[1945] = n_Body_x[1945];
                c_Body_y[1945] = n_Body_y[1945];
                c_Body_x[1946] = n_Body_x[1946];
                c_Body_y[1946] = n_Body_y[1946];
                c_Body_x[1947] = n_Body_x[1947];
                c_Body_y[1947] = n_Body_y[1947];
                c_Body_x[1948] = n_Body_x[1948];
                c_Body_y[1948] = n_Body_y[1948];
                c_Body_x[1949] = n_Body_x[1949];
                c_Body_y[1949] = n_Body_y[1949];
                c_Body_x[1950] = n_Body_x[1950];
                c_Body_y[1950] = n_Body_y[1950];
                c_Body_x[1951] = n_Body_x[1951];
                c_Body_y[1951] = n_Body_y[1951];
                c_Body_x[1952] = n_Body_x[1952];
                c_Body_y[1952] = n_Body_y[1952];
                c_Body_x[1953] = n_Body_x[1953];
                c_Body_y[1953] = n_Body_y[1953];
                c_Body_x[1954] = n_Body_x[1954];
                c_Body_y[1954] = n_Body_y[1954];
                c_Body_x[1955] = n_Body_x[1955];
                c_Body_y[1955] = n_Body_y[1955];
                c_Body_x[1956] = n_Body_x[1956];
                c_Body_y[1956] = n_Body_y[1956];
                c_Body_x[1957] = n_Body_x[1957];
                c_Body_y[1957] = n_Body_y[1957];
                c_Body_x[1958] = n_Body_x[1958];
                c_Body_y[1958] = n_Body_y[1958];
                c_Body_x[1959] = n_Body_x[1959];
                c_Body_y[1959] = n_Body_y[1959];
                c_Body_x[1960] = n_Body_x[1960];
                c_Body_y[1960] = n_Body_y[1960];
                c_Body_x[1961] = n_Body_x[1961];
                c_Body_y[1961] = n_Body_y[1961];
                c_Body_x[1962] = n_Body_x[1962];
                c_Body_y[1962] = n_Body_y[1962];
                c_Body_x[1963] = n_Body_x[1963];
                c_Body_y[1963] = n_Body_y[1963];
                c_Body_x[1964] = n_Body_x[1964];
                c_Body_y[1964] = n_Body_y[1964];
                c_Body_x[1965] = n_Body_x[1965];
                c_Body_y[1965] = n_Body_y[1965];
                c_Body_x[1966] = n_Body_x[1966];
                c_Body_y[1966] = n_Body_y[1966];
                c_Body_x[1967] = n_Body_x[1967];
                c_Body_y[1967] = n_Body_y[1967];
                c_Body_x[1968] = n_Body_x[1968];
                c_Body_y[1968] = n_Body_y[1968];
                c_Body_x[1969] = n_Body_x[1969];
                c_Body_y[1969] = n_Body_y[1969];
                c_Body_x[1970] = n_Body_x[1970];
                c_Body_y[1970] = n_Body_y[1970];
                c_Body_x[1971] = n_Body_x[1971];
                c_Body_y[1971] = n_Body_y[1971];
                c_Body_x[1972] = n_Body_x[1972];
                c_Body_y[1972] = n_Body_y[1972];
                c_Body_x[1973] = n_Body_x[1973];
                c_Body_y[1973] = n_Body_y[1973];
                c_Body_x[1974] = n_Body_x[1974];
                c_Body_y[1974] = n_Body_y[1974];
                c_Body_x[1975] = n_Body_x[1975];
                c_Body_y[1975] = n_Body_y[1975];
                c_Body_x[1976] = n_Body_x[1976];
                c_Body_y[1976] = n_Body_y[1976];
                c_Body_x[1977] = n_Body_x[1977];
                c_Body_y[1977] = n_Body_y[1977];
                c_Body_x[1978] = n_Body_x[1978];
                c_Body_y[1978] = n_Body_y[1978];
                c_Body_x[1979] = n_Body_x[1979];
                c_Body_y[1979] = n_Body_y[1979];
                c_Body_x[1980] = n_Body_x[1980];
                c_Body_y[1980] = n_Body_y[1980];
                c_Body_x[1981] = n_Body_x[1981];
                c_Body_y[1981] = n_Body_y[1981];
                c_Body_x[1982] = n_Body_x[1982];
                c_Body_y[1982] = n_Body_y[1982];
                c_Body_x[1983] = n_Body_x[1983];
                c_Body_y[1983] = n_Body_y[1983];
                c_Body_x[1984] = n_Body_x[1984];
                c_Body_y[1984] = n_Body_y[1984];
                c_Body_x[1985] = n_Body_x[1985];
                c_Body_y[1985] = n_Body_y[1985];
                c_Body_x[1986] = n_Body_x[1986];
                c_Body_y[1986] = n_Body_y[1986];
                c_Body_x[1987] = n_Body_x[1987];
                c_Body_y[1987] = n_Body_y[1987];
                c_Body_x[1988] = n_Body_x[1988];
                c_Body_y[1988] = n_Body_y[1988];
                c_Body_x[1989] = n_Body_x[1989];
                c_Body_y[1989] = n_Body_y[1989];
                c_Body_x[1990] = n_Body_x[1990];
                c_Body_y[1990] = n_Body_y[1990];
                c_Body_x[1991] = n_Body_x[1991];
                c_Body_y[1991] = n_Body_y[1991];
                c_Body_x[1992] = n_Body_x[1992];
                c_Body_y[1992] = n_Body_y[1992];
                c_Body_x[1993] = n_Body_x[1993];
                c_Body_y[1993] = n_Body_y[1993];
                c_Body_x[1994] = n_Body_x[1994];
                c_Body_y[1994] = n_Body_y[1994];
                c_Body_x[1995] = n_Body_x[1995];
                c_Body_y[1995] = n_Body_y[1995];
                c_Body_x[1996] = n_Body_x[1996];
                c_Body_y[1996] = n_Body_y[1996];
                c_Body_x[1997] = n_Body_x[1997];
                c_Body_y[1997] = n_Body_y[1997];
                c_Body_x[1998] = n_Body_x[1998];
                c_Body_y[1998] = n_Body_y[1998];
                c_Body_x[1999] = n_Body_x[1999];
                c_Body_y[1999] = n_Body_y[1999];
                c_Body_x[2000] = n_Body_x[2000];
                c_Body_y[2000] = n_Body_y[2000];
                c_Body_x[2001] = n_Body_x[2001];
                c_Body_y[2001] = n_Body_y[2001];
                c_Body_x[2002] = n_Body_x[2002];
                c_Body_y[2002] = n_Body_y[2002];
                c_Body_x[2003] = n_Body_x[2003];
                c_Body_y[2003] = n_Body_y[2003];
                c_Body_x[2004] = n_Body_x[2004];
                c_Body_y[2004] = n_Body_y[2004];
                c_Body_x[2005] = n_Body_x[2005];
                c_Body_y[2005] = n_Body_y[2005];
                c_Body_x[2006] = n_Body_x[2006];
                c_Body_y[2006] = n_Body_y[2006];
                c_Body_x[2007] = n_Body_x[2007];
                c_Body_y[2007] = n_Body_y[2007];
                c_Body_x[2008] = n_Body_x[2008];
                c_Body_y[2008] = n_Body_y[2008];
                c_Body_x[2009] = n_Body_x[2009];
                c_Body_y[2009] = n_Body_y[2009];
                c_Body_x[2010] = n_Body_x[2010];
                c_Body_y[2010] = n_Body_y[2010];
                c_Body_x[2011] = n_Body_x[2011];
                c_Body_y[2011] = n_Body_y[2011];
                c_Body_x[2012] = n_Body_x[2012];
                c_Body_y[2012] = n_Body_y[2012];
                c_Body_x[2013] = n_Body_x[2013];
                c_Body_y[2013] = n_Body_y[2013];
                c_Body_x[2014] = n_Body_x[2014];
                c_Body_y[2014] = n_Body_y[2014];
                c_Body_x[2015] = n_Body_x[2015];
                c_Body_y[2015] = n_Body_y[2015];
                c_Body_x[2016] = n_Body_x[2016];
                c_Body_y[2016] = n_Body_y[2016];
                c_Body_x[2017] = n_Body_x[2017];
                c_Body_y[2017] = n_Body_y[2017];
                c_Body_x[2018] = n_Body_x[2018];
                c_Body_y[2018] = n_Body_y[2018];
                c_Body_x[2019] = n_Body_x[2019];
                c_Body_y[2019] = n_Body_y[2019];
                c_Body_x[2020] = n_Body_x[2020];
                c_Body_y[2020] = n_Body_y[2020];
                c_Body_x[2021] = n_Body_x[2021];
                c_Body_y[2021] = n_Body_y[2021];
                c_Body_x[2022] = n_Body_x[2022];
                c_Body_y[2022] = n_Body_y[2022];
                c_Body_x[2023] = n_Body_x[2023];
                c_Body_y[2023] = n_Body_y[2023];
                c_Body_x[2024] = n_Body_x[2024];
                c_Body_y[2024] = n_Body_y[2024];
                c_Body_x[2025] = n_Body_x[2025];
                c_Body_y[2025] = n_Body_y[2025];
                c_Body_x[2026] = n_Body_x[2026];
                c_Body_y[2026] = n_Body_y[2026];
                c_Body_x[2027] = n_Body_x[2027];
                c_Body_y[2027] = n_Body_y[2027];
                c_Body_x[2028] = n_Body_x[2028];
                c_Body_y[2028] = n_Body_y[2028];
                c_Body_x[2029] = n_Body_x[2029];
                c_Body_y[2029] = n_Body_y[2029];
                c_Body_x[2030] = n_Body_x[2030];
                c_Body_y[2030] = n_Body_y[2030];
                c_Body_x[2031] = n_Body_x[2031];
                c_Body_y[2031] = n_Body_y[2031];
                c_Body_x[2032] = n_Body_x[2032];
                c_Body_y[2032] = n_Body_y[2032];
                c_Body_x[2033] = n_Body_x[2033];
                c_Body_y[2033] = n_Body_y[2033];
                c_Body_x[2034] = n_Body_x[2034];
                c_Body_y[2034] = n_Body_y[2034];
                c_Body_x[2035] = n_Body_x[2035];
                c_Body_y[2035] = n_Body_y[2035];
                c_Body_x[2036] = n_Body_x[2036];
                c_Body_y[2036] = n_Body_y[2036];
                c_Body_x[2037] = n_Body_x[2037];
                c_Body_y[2037] = n_Body_y[2037];
                c_Body_x[2038] = n_Body_x[2038];
                c_Body_y[2038] = n_Body_y[2038];
                c_Body_x[2039] = n_Body_x[2039];
                c_Body_y[2039] = n_Body_y[2039];
                c_Body_x[2040] = n_Body_x[2040];
                c_Body_y[2040] = n_Body_y[2040];
                c_Body_x[2041] = n_Body_x[2041];
                c_Body_y[2041] = n_Body_y[2041];
                c_Body_x[2042] = n_Body_x[2042];
                c_Body_y[2042] = n_Body_y[2042];
                c_Body_x[2043] = n_Body_x[2043];
                c_Body_y[2043] = n_Body_y[2043];
                c_Body_x[2044] = n_Body_x[2044];
                c_Body_y[2044] = n_Body_y[2044];
                c_Body_x[2045] = n_Body_x[2045];
                c_Body_y[2045] = n_Body_y[2045];
                c_Body_x[2046] = n_Body_x[2046];
                c_Body_y[2046] = n_Body_y[2046];
                c_Body_x[2047] = n_Body_x[2047];
                c_Body_y[2047] = n_Body_y[2047];
                c_Body_x[2048] = n_Body_x[2048];
                c_Body_y[2048] = n_Body_y[2048];
                c_Body_x[2049] = n_Body_x[2049];
                c_Body_y[2049] = n_Body_y[2049];
                c_Body_x[2050] = n_Body_x[2050];
                c_Body_y[2050] = n_Body_y[2050];
                c_Body_x[2051] = n_Body_x[2051];
                c_Body_y[2051] = n_Body_y[2051];
                c_Body_x[2052] = n_Body_x[2052];
                c_Body_y[2052] = n_Body_y[2052];
                c_Body_x[2053] = n_Body_x[2053];
                c_Body_y[2053] = n_Body_y[2053];
                c_Body_x[2054] = n_Body_x[2054];
                c_Body_y[2054] = n_Body_y[2054];
                c_Body_x[2055] = n_Body_x[2055];
                c_Body_y[2055] = n_Body_y[2055];
                c_Body_x[2056] = n_Body_x[2056];
                c_Body_y[2056] = n_Body_y[2056];
                c_Body_x[2057] = n_Body_x[2057];
                c_Body_y[2057] = n_Body_y[2057];
                c_Body_x[2058] = n_Body_x[2058];
                c_Body_y[2058] = n_Body_y[2058];
                c_Body_x[2059] = n_Body_x[2059];
                c_Body_y[2059] = n_Body_y[2059];
                c_Body_x[2060] = n_Body_x[2060];
                c_Body_y[2060] = n_Body_y[2060];
                c_Body_x[2061] = n_Body_x[2061];
                c_Body_y[2061] = n_Body_y[2061];
                c_Body_x[2062] = n_Body_x[2062];
                c_Body_y[2062] = n_Body_y[2062];
                c_Body_x[2063] = n_Body_x[2063];
                c_Body_y[2063] = n_Body_y[2063];
                c_Body_x[2064] = n_Body_x[2064];
                c_Body_y[2064] = n_Body_y[2064];
                c_Body_x[2065] = n_Body_x[2065];
                c_Body_y[2065] = n_Body_y[2065];
                c_Body_x[2066] = n_Body_x[2066];
                c_Body_y[2066] = n_Body_y[2066];
                c_Body_x[2067] = n_Body_x[2067];
                c_Body_y[2067] = n_Body_y[2067];
                c_Body_x[2068] = n_Body_x[2068];
                c_Body_y[2068] = n_Body_y[2068];
                c_Body_x[2069] = n_Body_x[2069];
                c_Body_y[2069] = n_Body_y[2069];
                c_Body_x[2070] = n_Body_x[2070];
                c_Body_y[2070] = n_Body_y[2070];
                c_Body_x[2071] = n_Body_x[2071];
                c_Body_y[2071] = n_Body_y[2071];
                c_Body_x[2072] = n_Body_x[2072];
                c_Body_y[2072] = n_Body_y[2072];
                c_Body_x[2073] = n_Body_x[2073];
                c_Body_y[2073] = n_Body_y[2073];
                c_Body_x[2074] = n_Body_x[2074];
                c_Body_y[2074] = n_Body_y[2074];
                c_Body_x[2075] = n_Body_x[2075];
                c_Body_y[2075] = n_Body_y[2075];
                c_Body_x[2076] = n_Body_x[2076];
                c_Body_y[2076] = n_Body_y[2076];
                c_Body_x[2077] = n_Body_x[2077];
                c_Body_y[2077] = n_Body_y[2077];
                c_Body_x[2078] = n_Body_x[2078];
                c_Body_y[2078] = n_Body_y[2078];
                c_Body_x[2079] = n_Body_x[2079];
                c_Body_y[2079] = n_Body_y[2079];
                c_Body_x[2080] = n_Body_x[2080];
                c_Body_y[2080] = n_Body_y[2080];
                c_Body_x[2081] = n_Body_x[2081];
                c_Body_y[2081] = n_Body_y[2081];
                c_Body_x[2082] = n_Body_x[2082];
                c_Body_y[2082] = n_Body_y[2082];
                c_Body_x[2083] = n_Body_x[2083];
                c_Body_y[2083] = n_Body_y[2083];
                c_Body_x[2084] = n_Body_x[2084];
                c_Body_y[2084] = n_Body_y[2084];
                c_Body_x[2085] = n_Body_x[2085];
                c_Body_y[2085] = n_Body_y[2085];
                c_Body_x[2086] = n_Body_x[2086];
                c_Body_y[2086] = n_Body_y[2086];
                c_Body_x[2087] = n_Body_x[2087];
                c_Body_y[2087] = n_Body_y[2087];
                c_Body_x[2088] = n_Body_x[2088];
                c_Body_y[2088] = n_Body_y[2088];
                c_Body_x[2089] = n_Body_x[2089];
                c_Body_y[2089] = n_Body_y[2089];
                c_Body_x[2090] = n_Body_x[2090];
                c_Body_y[2090] = n_Body_y[2090];
                c_Body_x[2091] = n_Body_x[2091];
                c_Body_y[2091] = n_Body_y[2091];
                c_Body_x[2092] = n_Body_x[2092];
                c_Body_y[2092] = n_Body_y[2092];
                c_Body_x[2093] = n_Body_x[2093];
                c_Body_y[2093] = n_Body_y[2093];
                c_Body_x[2094] = n_Body_x[2094];
                c_Body_y[2094] = n_Body_y[2094];
                c_Body_x[2095] = n_Body_x[2095];
                c_Body_y[2095] = n_Body_y[2095];
                c_Body_x[2096] = n_Body_x[2096];
                c_Body_y[2096] = n_Body_y[2096];
                c_Body_x[2097] = n_Body_x[2097];
                c_Body_y[2097] = n_Body_y[2097];
                c_Body_x[2098] = n_Body_x[2098];
                c_Body_y[2098] = n_Body_y[2098];
                c_Body_x[2099] = n_Body_x[2099];
                c_Body_y[2099] = n_Body_y[2099];
                c_Body_x[2100] = n_Body_x[2100];
                c_Body_y[2100] = n_Body_y[2100];
                c_Body_x[2101] = n_Body_x[2101];
                c_Body_y[2101] = n_Body_y[2101];
                c_Body_x[2102] = n_Body_x[2102];
                c_Body_y[2102] = n_Body_y[2102];
                c_Body_x[2103] = n_Body_x[2103];
                c_Body_y[2103] = n_Body_y[2103];
                c_Body_x[2104] = n_Body_x[2104];
                c_Body_y[2104] = n_Body_y[2104];
                c_Body_x[2105] = n_Body_x[2105];
                c_Body_y[2105] = n_Body_y[2105];
                c_Body_x[2106] = n_Body_x[2106];
                c_Body_y[2106] = n_Body_y[2106];
                c_Body_x[2107] = n_Body_x[2107];
                c_Body_y[2107] = n_Body_y[2107];
                c_Body_x[2108] = n_Body_x[2108];
                c_Body_y[2108] = n_Body_y[2108];
                c_Body_x[2109] = n_Body_x[2109];
                c_Body_y[2109] = n_Body_y[2109];
                c_Body_x[2110] = n_Body_x[2110];
                c_Body_y[2110] = n_Body_y[2110];
                c_Body_x[2111] = n_Body_x[2111];
                c_Body_y[2111] = n_Body_y[2111];
                c_Body_x[2112] = n_Body_x[2112];
                c_Body_y[2112] = n_Body_y[2112];
                c_Body_x[2113] = n_Body_x[2113];
                c_Body_y[2113] = n_Body_y[2113];
                c_Body_x[2114] = n_Body_x[2114];
                c_Body_y[2114] = n_Body_y[2114];
                c_Body_x[2115] = n_Body_x[2115];
                c_Body_y[2115] = n_Body_y[2115];
                c_Body_x[2116] = n_Body_x[2116];
                c_Body_y[2116] = n_Body_y[2116];
                c_Body_x[2117] = n_Body_x[2117];
                c_Body_y[2117] = n_Body_y[2117];
                c_Body_x[2118] = n_Body_x[2118];
                c_Body_y[2118] = n_Body_y[2118];
                c_Body_x[2119] = n_Body_x[2119];
                c_Body_y[2119] = n_Body_y[2119];
                c_Body_x[2120] = n_Body_x[2120];
                c_Body_y[2120] = n_Body_y[2120];
                c_Body_x[2121] = n_Body_x[2121];
                c_Body_y[2121] = n_Body_y[2121];
                c_Body_x[2122] = n_Body_x[2122];
                c_Body_y[2122] = n_Body_y[2122];
                c_Body_x[2123] = n_Body_x[2123];
                c_Body_y[2123] = n_Body_y[2123];
                c_Body_x[2124] = n_Body_x[2124];
                c_Body_y[2124] = n_Body_y[2124];
                c_Body_x[2125] = n_Body_x[2125];
                c_Body_y[2125] = n_Body_y[2125];
                c_Body_x[2126] = n_Body_x[2126];
                c_Body_y[2126] = n_Body_y[2126];
                c_Body_x[2127] = n_Body_x[2127];
                c_Body_y[2127] = n_Body_y[2127];
                c_Body_x[2128] = n_Body_x[2128];
                c_Body_y[2128] = n_Body_y[2128];
                c_Body_x[2129] = n_Body_x[2129];
                c_Body_y[2129] = n_Body_y[2129];
                c_Body_x[2130] = n_Body_x[2130];
                c_Body_y[2130] = n_Body_y[2130];
                c_Body_x[2131] = n_Body_x[2131];
                c_Body_y[2131] = n_Body_y[2131];
                c_Body_x[2132] = n_Body_x[2132];
                c_Body_y[2132] = n_Body_y[2132];
                c_Body_x[2133] = n_Body_x[2133];
                c_Body_y[2133] = n_Body_y[2133];
                c_Body_x[2134] = n_Body_x[2134];
                c_Body_y[2134] = n_Body_y[2134];
                c_Body_x[2135] = n_Body_x[2135];
                c_Body_y[2135] = n_Body_y[2135];
                c_Body_x[2136] = n_Body_x[2136];
                c_Body_y[2136] = n_Body_y[2136];
                c_Body_x[2137] = n_Body_x[2137];
                c_Body_y[2137] = n_Body_y[2137];
                c_Body_x[2138] = n_Body_x[2138];
                c_Body_y[2138] = n_Body_y[2138];
                c_Body_x[2139] = n_Body_x[2139];
                c_Body_y[2139] = n_Body_y[2139];
                c_Body_x[2140] = n_Body_x[2140];
                c_Body_y[2140] = n_Body_y[2140];
                c_Body_x[2141] = n_Body_x[2141];
                c_Body_y[2141] = n_Body_y[2141];
                c_Body_x[2142] = n_Body_x[2142];
                c_Body_y[2142] = n_Body_y[2142];
                c_Body_x[2143] = n_Body_x[2143];
                c_Body_y[2143] = n_Body_y[2143];
                c_Body_x[2144] = n_Body_x[2144];
                c_Body_y[2144] = n_Body_y[2144];
                c_Body_x[2145] = n_Body_x[2145];
                c_Body_y[2145] = n_Body_y[2145];
                c_Body_x[2146] = n_Body_x[2146];
                c_Body_y[2146] = n_Body_y[2146];
                c_Body_x[2147] = n_Body_x[2147];
                c_Body_y[2147] = n_Body_y[2147];
                c_Body_x[2148] = n_Body_x[2148];
                c_Body_y[2148] = n_Body_y[2148];
                c_Body_x[2149] = n_Body_x[2149];
                c_Body_y[2149] = n_Body_y[2149];
                c_Body_x[2150] = n_Body_x[2150];
                c_Body_y[2150] = n_Body_y[2150];
                c_Body_x[2151] = n_Body_x[2151];
                c_Body_y[2151] = n_Body_y[2151];
                c_Body_x[2152] = n_Body_x[2152];
                c_Body_y[2152] = n_Body_y[2152];
                c_Body_x[2153] = n_Body_x[2153];
                c_Body_y[2153] = n_Body_y[2153];
                c_Body_x[2154] = n_Body_x[2154];
                c_Body_y[2154] = n_Body_y[2154];
                c_Body_x[2155] = n_Body_x[2155];
                c_Body_y[2155] = n_Body_y[2155];
                c_Body_x[2156] = n_Body_x[2156];
                c_Body_y[2156] = n_Body_y[2156];
                c_Body_x[2157] = n_Body_x[2157];
                c_Body_y[2157] = n_Body_y[2157];
                c_Body_x[2158] = n_Body_x[2158];
                c_Body_y[2158] = n_Body_y[2158];
                c_Body_x[2159] = n_Body_x[2159];
                c_Body_y[2159] = n_Body_y[2159];
                c_Body_x[2160] = n_Body_x[2160];
                c_Body_y[2160] = n_Body_y[2160];
                c_Body_x[2161] = n_Body_x[2161];
                c_Body_y[2161] = n_Body_y[2161];
                c_Body_x[2162] = n_Body_x[2162];
                c_Body_y[2162] = n_Body_y[2162];
                c_Body_x[2163] = n_Body_x[2163];
                c_Body_y[2163] = n_Body_y[2163];
                c_Body_x[2164] = n_Body_x[2164];
                c_Body_y[2164] = n_Body_y[2164];
                c_Body_x[2165] = n_Body_x[2165];
                c_Body_y[2165] = n_Body_y[2165];
                c_Body_x[2166] = n_Body_x[2166];
                c_Body_y[2166] = n_Body_y[2166];
                c_Body_x[2167] = n_Body_x[2167];
                c_Body_y[2167] = n_Body_y[2167];
                c_Body_x[2168] = n_Body_x[2168];
                c_Body_y[2168] = n_Body_y[2168];
                c_Body_x[2169] = n_Body_x[2169];
                c_Body_y[2169] = n_Body_y[2169];
                c_Body_x[2170] = n_Body_x[2170];
                c_Body_y[2170] = n_Body_y[2170];
                c_Body_x[2171] = n_Body_x[2171];
                c_Body_y[2171] = n_Body_y[2171];
                c_Body_x[2172] = n_Body_x[2172];
                c_Body_y[2172] = n_Body_y[2172];
                c_Body_x[2173] = n_Body_x[2173];
                c_Body_y[2173] = n_Body_y[2173];
                c_Body_x[2174] = n_Body_x[2174];
                c_Body_y[2174] = n_Body_y[2174];
                c_Body_x[2175] = n_Body_x[2175];
                c_Body_y[2175] = n_Body_y[2175];
                c_Body_x[2176] = n_Body_x[2176];
                c_Body_y[2176] = n_Body_y[2176];
                c_Body_x[2177] = n_Body_x[2177];
                c_Body_y[2177] = n_Body_y[2177];
                c_Body_x[2178] = n_Body_x[2178];
                c_Body_y[2178] = n_Body_y[2178];
                c_Body_x[2179] = n_Body_x[2179];
                c_Body_y[2179] = n_Body_y[2179];
                c_Body_x[2180] = n_Body_x[2180];
                c_Body_y[2180] = n_Body_y[2180];
                c_Body_x[2181] = n_Body_x[2181];
                c_Body_y[2181] = n_Body_y[2181];
                c_Body_x[2182] = n_Body_x[2182];
                c_Body_y[2182] = n_Body_y[2182];
                c_Body_x[2183] = n_Body_x[2183];
                c_Body_y[2183] = n_Body_y[2183];
                c_Body_x[2184] = n_Body_x[2184];
                c_Body_y[2184] = n_Body_y[2184];
                c_Body_x[2185] = n_Body_x[2185];
                c_Body_y[2185] = n_Body_y[2185];
                c_Body_x[2186] = n_Body_x[2186];
                c_Body_y[2186] = n_Body_y[2186];
                c_Body_x[2187] = n_Body_x[2187];
                c_Body_y[2187] = n_Body_y[2187];
                c_Body_x[2188] = n_Body_x[2188];
                c_Body_y[2188] = n_Body_y[2188];
                c_Body_x[2189] = n_Body_x[2189];
                c_Body_y[2189] = n_Body_y[2189];
                c_Body_x[2190] = n_Body_x[2190];
                c_Body_y[2190] = n_Body_y[2190];
                c_Body_x[2191] = n_Body_x[2191];
                c_Body_y[2191] = n_Body_y[2191];
                c_Body_x[2192] = n_Body_x[2192];
                c_Body_y[2192] = n_Body_y[2192];
                c_Body_x[2193] = n_Body_x[2193];
                c_Body_y[2193] = n_Body_y[2193];
                c_Body_x[2194] = n_Body_x[2194];
                c_Body_y[2194] = n_Body_y[2194];
                c_Body_x[2195] = n_Body_x[2195];
                c_Body_y[2195] = n_Body_y[2195];
                c_Body_x[2196] = n_Body_x[2196];
                c_Body_y[2196] = n_Body_y[2196];
                c_Body_x[2197] = n_Body_x[2197];
                c_Body_y[2197] = n_Body_y[2197];
                c_Body_x[2198] = n_Body_x[2198];
                c_Body_y[2198] = n_Body_y[2198];
                c_Body_x[2199] = n_Body_x[2199];
                c_Body_y[2199] = n_Body_y[2199];
                c_Body_x[2200] = n_Body_x[2200];
                c_Body_y[2200] = n_Body_y[2200];
                c_Body_x[2201] = n_Body_x[2201];
                c_Body_y[2201] = n_Body_y[2201];
                c_Body_x[2202] = n_Body_x[2202];
                c_Body_y[2202] = n_Body_y[2202];
                c_Body_x[2203] = n_Body_x[2203];
                c_Body_y[2203] = n_Body_y[2203];
                c_Body_x[2204] = n_Body_x[2204];
                c_Body_y[2204] = n_Body_y[2204];
                c_Body_x[2205] = n_Body_x[2205];
                c_Body_y[2205] = n_Body_y[2205];
                c_Body_x[2206] = n_Body_x[2206];
                c_Body_y[2206] = n_Body_y[2206];
                c_Body_x[2207] = n_Body_x[2207];
                c_Body_y[2207] = n_Body_y[2207];
                c_Body_x[2208] = n_Body_x[2208];
                c_Body_y[2208] = n_Body_y[2208];
                c_Body_x[2209] = n_Body_x[2209];
                c_Body_y[2209] = n_Body_y[2209];
                c_Body_x[2210] = n_Body_x[2210];
                c_Body_y[2210] = n_Body_y[2210];
                c_Body_x[2211] = n_Body_x[2211];
                c_Body_y[2211] = n_Body_y[2211];
                c_Body_x[2212] = n_Body_x[2212];
                c_Body_y[2212] = n_Body_y[2212];
                c_Body_x[2213] = n_Body_x[2213];
                c_Body_y[2213] = n_Body_y[2213];
                c_Body_x[2214] = n_Body_x[2214];
                c_Body_y[2214] = n_Body_y[2214];
                c_Body_x[2215] = n_Body_x[2215];
                c_Body_y[2215] = n_Body_y[2215];
                c_Body_x[2216] = n_Body_x[2216];
                c_Body_y[2216] = n_Body_y[2216];
                c_Body_x[2217] = n_Body_x[2217];
                c_Body_y[2217] = n_Body_y[2217];
                c_Body_x[2218] = n_Body_x[2218];
                c_Body_y[2218] = n_Body_y[2218];
                c_Body_x[2219] = n_Body_x[2219];
                c_Body_y[2219] = n_Body_y[2219];
                c_Body_x[2220] = n_Body_x[2220];
                c_Body_y[2220] = n_Body_y[2220];
                c_Body_x[2221] = n_Body_x[2221];
                c_Body_y[2221] = n_Body_y[2221];
                c_Body_x[2222] = n_Body_x[2222];
                c_Body_y[2222] = n_Body_y[2222];
                c_Body_x[2223] = n_Body_x[2223];
                c_Body_y[2223] = n_Body_y[2223];
                c_Body_x[2224] = n_Body_x[2224];
                c_Body_y[2224] = n_Body_y[2224];
                c_Body_x[2225] = n_Body_x[2225];
                c_Body_y[2225] = n_Body_y[2225];
                c_Body_x[2226] = n_Body_x[2226];
                c_Body_y[2226] = n_Body_y[2226];
                c_Body_x[2227] = n_Body_x[2227];
                c_Body_y[2227] = n_Body_y[2227];
                c_Body_x[2228] = n_Body_x[2228];
                c_Body_y[2228] = n_Body_y[2228];
                c_Body_x[2229] = n_Body_x[2229];
                c_Body_y[2229] = n_Body_y[2229];
                c_Body_x[2230] = n_Body_x[2230];
                c_Body_y[2230] = n_Body_y[2230];
                c_Body_x[2231] = n_Body_x[2231];
                c_Body_y[2231] = n_Body_y[2231];
                c_Body_x[2232] = n_Body_x[2232];
                c_Body_y[2232] = n_Body_y[2232];
                c_Body_x[2233] = n_Body_x[2233];
                c_Body_y[2233] = n_Body_y[2233];
                c_Body_x[2234] = n_Body_x[2234];
                c_Body_y[2234] = n_Body_y[2234];
                c_Body_x[2235] = n_Body_x[2235];
                c_Body_y[2235] = n_Body_y[2235];
                c_Body_x[2236] = n_Body_x[2236];
                c_Body_y[2236] = n_Body_y[2236];
                c_Body_x[2237] = n_Body_x[2237];
                c_Body_y[2237] = n_Body_y[2237];
                c_Body_x[2238] = n_Body_x[2238];
                c_Body_y[2238] = n_Body_y[2238];
                c_Body_x[2239] = n_Body_x[2239];
                c_Body_y[2239] = n_Body_y[2239];
                c_Body_x[2240] = n_Body_x[2240];
                c_Body_y[2240] = n_Body_y[2240];
                c_Body_x[2241] = n_Body_x[2241];
                c_Body_y[2241] = n_Body_y[2241];
                c_Body_x[2242] = n_Body_x[2242];
                c_Body_y[2242] = n_Body_y[2242];
                c_Body_x[2243] = n_Body_x[2243];
                c_Body_y[2243] = n_Body_y[2243];
                c_Body_x[2244] = n_Body_x[2244];
                c_Body_y[2244] = n_Body_y[2244];
                c_Body_x[2245] = n_Body_x[2245];
                c_Body_y[2245] = n_Body_y[2245];
                c_Body_x[2246] = n_Body_x[2246];
                c_Body_y[2246] = n_Body_y[2246];
                c_Body_x[2247] = n_Body_x[2247];
                c_Body_y[2247] = n_Body_y[2247];
                c_Body_x[2248] = n_Body_x[2248];
                c_Body_y[2248] = n_Body_y[2248];
                c_Body_x[2249] = n_Body_x[2249];
                c_Body_y[2249] = n_Body_y[2249];
                c_Body_x[2250] = n_Body_x[2250];
                c_Body_y[2250] = n_Body_y[2250];
                c_Body_x[2251] = n_Body_x[2251];
                c_Body_y[2251] = n_Body_y[2251];
                c_Body_x[2252] = n_Body_x[2252];
                c_Body_y[2252] = n_Body_y[2252];
                c_Body_x[2253] = n_Body_x[2253];
                c_Body_y[2253] = n_Body_y[2253];
                c_Body_x[2254] = n_Body_x[2254];
                c_Body_y[2254] = n_Body_y[2254];
                c_Body_x[2255] = n_Body_x[2255];
                c_Body_y[2255] = n_Body_y[2255];
                c_Body_x[2256] = n_Body_x[2256];
                c_Body_y[2256] = n_Body_y[2256];
                c_Body_x[2257] = n_Body_x[2257];
                c_Body_y[2257] = n_Body_y[2257];
                c_Body_x[2258] = n_Body_x[2258];
                c_Body_y[2258] = n_Body_y[2258];
                c_Body_x[2259] = n_Body_x[2259];
                c_Body_y[2259] = n_Body_y[2259];
                c_Body_x[2260] = n_Body_x[2260];
                c_Body_y[2260] = n_Body_y[2260];
                c_Body_x[2261] = n_Body_x[2261];
                c_Body_y[2261] = n_Body_y[2261];
                c_Body_x[2262] = n_Body_x[2262];
                c_Body_y[2262] = n_Body_y[2262];
                c_Body_x[2263] = n_Body_x[2263];
                c_Body_y[2263] = n_Body_y[2263];
                c_Body_x[2264] = n_Body_x[2264];
                c_Body_y[2264] = n_Body_y[2264];
                c_Body_x[2265] = n_Body_x[2265];
                c_Body_y[2265] = n_Body_y[2265];
                c_Body_x[2266] = n_Body_x[2266];
                c_Body_y[2266] = n_Body_y[2266];
                c_Body_x[2267] = n_Body_x[2267];
                c_Body_y[2267] = n_Body_y[2267];
                c_Body_x[2268] = n_Body_x[2268];
                c_Body_y[2268] = n_Body_y[2268];
                c_Body_x[2269] = n_Body_x[2269];
                c_Body_y[2269] = n_Body_y[2269];
                c_Body_x[2270] = n_Body_x[2270];
                c_Body_y[2270] = n_Body_y[2270];
                c_Body_x[2271] = n_Body_x[2271];
                c_Body_y[2271] = n_Body_y[2271];
                c_Body_x[2272] = n_Body_x[2272];
                c_Body_y[2272] = n_Body_y[2272];
                c_Body_x[2273] = n_Body_x[2273];
                c_Body_y[2273] = n_Body_y[2273];
                c_Body_x[2274] = n_Body_x[2274];
                c_Body_y[2274] = n_Body_y[2274];
                c_Body_x[2275] = n_Body_x[2275];
                c_Body_y[2275] = n_Body_y[2275];
                c_Body_x[2276] = n_Body_x[2276];
                c_Body_y[2276] = n_Body_y[2276];
                c_Body_x[2277] = n_Body_x[2277];
                c_Body_y[2277] = n_Body_y[2277];
                c_Body_x[2278] = n_Body_x[2278];
                c_Body_y[2278] = n_Body_y[2278];
                c_Body_x[2279] = n_Body_x[2279];
                c_Body_y[2279] = n_Body_y[2279];
                c_Body_x[2280] = n_Body_x[2280];
                c_Body_y[2280] = n_Body_y[2280];
                c_Body_x[2281] = n_Body_x[2281];
                c_Body_y[2281] = n_Body_y[2281];
                c_Body_x[2282] = n_Body_x[2282];
                c_Body_y[2282] = n_Body_y[2282];
                c_Body_x[2283] = n_Body_x[2283];
                c_Body_y[2283] = n_Body_y[2283];
                c_Body_x[2284] = n_Body_x[2284];
                c_Body_y[2284] = n_Body_y[2284];
                c_Body_x[2285] = n_Body_x[2285];
                c_Body_y[2285] = n_Body_y[2285];
                c_Body_x[2286] = n_Body_x[2286];
                c_Body_y[2286] = n_Body_y[2286];
                c_Body_x[2287] = n_Body_x[2287];
                c_Body_y[2287] = n_Body_y[2287];
                c_Body_x[2288] = n_Body_x[2288];
                c_Body_y[2288] = n_Body_y[2288];
                c_Body_x[2289] = n_Body_x[2289];
                c_Body_y[2289] = n_Body_y[2289];
                c_Body_x[2290] = n_Body_x[2290];
                c_Body_y[2290] = n_Body_y[2290];
                c_Body_x[2291] = n_Body_x[2291];
                c_Body_y[2291] = n_Body_y[2291];
                c_Body_x[2292] = n_Body_x[2292];
                c_Body_y[2292] = n_Body_y[2292];
                c_Body_x[2293] = n_Body_x[2293];
                c_Body_y[2293] = n_Body_y[2293];
                c_Body_x[2294] = n_Body_x[2294];
                c_Body_y[2294] = n_Body_y[2294];
                c_Body_x[2295] = n_Body_x[2295];
                c_Body_y[2295] = n_Body_y[2295];
                c_Body_x[2296] = n_Body_x[2296];
                c_Body_y[2296] = n_Body_y[2296];
                c_Body_x[2297] = n_Body_x[2297];
                c_Body_y[2297] = n_Body_y[2297];
                c_Body_x[2298] = n_Body_x[2298];
                c_Body_y[2298] = n_Body_y[2298];
                c_Body_x[2299] = n_Body_x[2299];
                c_Body_y[2299] = n_Body_y[2299];
                c_Body_x[2300] = n_Body_x[2300];
                c_Body_y[2300] = n_Body_y[2300];
                c_Body_x[2301] = n_Body_x[2301];
                c_Body_y[2301] = n_Body_y[2301];
                c_Body_x[2302] = n_Body_x[2302];
                c_Body_y[2302] = n_Body_y[2302];
                c_Body_x[2303] = n_Body_x[2303];
                c_Body_y[2303] = n_Body_y[2303];
                c_Body_x[2304] = n_Body_x[2304];
                c_Body_y[2304] = n_Body_y[2304];
                c_Body_x[2305] = n_Body_x[2305];
                c_Body_y[2305] = n_Body_y[2305];
                c_Body_x[2306] = n_Body_x[2306];
                c_Body_y[2306] = n_Body_y[2306];
                c_Body_x[2307] = n_Body_x[2307];
                c_Body_y[2307] = n_Body_y[2307];
                c_Body_x[2308] = n_Body_x[2308];
                c_Body_y[2308] = n_Body_y[2308];
                c_Body_x[2309] = n_Body_x[2309];
                c_Body_y[2309] = n_Body_y[2309];
                c_Body_x[2310] = n_Body_x[2310];
                c_Body_y[2310] = n_Body_y[2310];
                c_Body_x[2311] = n_Body_x[2311];
                c_Body_y[2311] = n_Body_y[2311];
                c_Body_x[2312] = n_Body_x[2312];
                c_Body_y[2312] = n_Body_y[2312];
                c_Body_x[2313] = n_Body_x[2313];
                c_Body_y[2313] = n_Body_y[2313];
                c_Body_x[2314] = n_Body_x[2314];
                c_Body_y[2314] = n_Body_y[2314];
                c_Body_x[2315] = n_Body_x[2315];
                c_Body_y[2315] = n_Body_y[2315];
                c_Body_x[2316] = n_Body_x[2316];
                c_Body_y[2316] = n_Body_y[2316];
                c_Body_x[2317] = n_Body_x[2317];
                c_Body_y[2317] = n_Body_y[2317];
                c_Body_x[2318] = n_Body_x[2318];
                c_Body_y[2318] = n_Body_y[2318];
                c_Body_x[2319] = n_Body_x[2319];
                c_Body_y[2319] = n_Body_y[2319];
                c_Body_x[2320] = n_Body_x[2320];
                c_Body_y[2320] = n_Body_y[2320];
                c_Body_x[2321] = n_Body_x[2321];
                c_Body_y[2321] = n_Body_y[2321];
                c_Body_x[2322] = n_Body_x[2322];
                c_Body_y[2322] = n_Body_y[2322];
                c_Body_x[2323] = n_Body_x[2323];
                c_Body_y[2323] = n_Body_y[2323];
                c_Body_x[2324] = n_Body_x[2324];
                c_Body_y[2324] = n_Body_y[2324];
                c_Body_x[2325] = n_Body_x[2325];
                c_Body_y[2325] = n_Body_y[2325];
                c_Body_x[2326] = n_Body_x[2326];
                c_Body_y[2326] = n_Body_y[2326];
                c_Body_x[2327] = n_Body_x[2327];
                c_Body_y[2327] = n_Body_y[2327];
                c_Body_x[2328] = n_Body_x[2328];
                c_Body_y[2328] = n_Body_y[2328];
                c_Body_x[2329] = n_Body_x[2329];
                c_Body_y[2329] = n_Body_y[2329];
                c_Body_x[2330] = n_Body_x[2330];
                c_Body_y[2330] = n_Body_y[2330];
                c_Body_x[2331] = n_Body_x[2331];
                c_Body_y[2331] = n_Body_y[2331];
                c_Body_x[2332] = n_Body_x[2332];
                c_Body_y[2332] = n_Body_y[2332];
                c_Body_x[2333] = n_Body_x[2333];
                c_Body_y[2333] = n_Body_y[2333];
                c_Body_x[2334] = n_Body_x[2334];
                c_Body_y[2334] = n_Body_y[2334];
                c_Body_x[2335] = n_Body_x[2335];
                c_Body_y[2335] = n_Body_y[2335];
                c_Body_x[2336] = n_Body_x[2336];
                c_Body_y[2336] = n_Body_y[2336];
                c_Body_x[2337] = n_Body_x[2337];
                c_Body_y[2337] = n_Body_y[2337];
                c_Body_x[2338] = n_Body_x[2338];
                c_Body_y[2338] = n_Body_y[2338];
                c_Body_x[2339] = n_Body_x[2339];
                c_Body_y[2339] = n_Body_y[2339];
                c_Body_x[2340] = n_Body_x[2340];
                c_Body_y[2340] = n_Body_y[2340];
                c_Body_x[2341] = n_Body_x[2341];
                c_Body_y[2341] = n_Body_y[2341];
                c_Body_x[2342] = n_Body_x[2342];
                c_Body_y[2342] = n_Body_y[2342];
                c_Body_x[2343] = n_Body_x[2343];
                c_Body_y[2343] = n_Body_y[2343];
                c_Body_x[2344] = n_Body_x[2344];
                c_Body_y[2344] = n_Body_y[2344];
                c_Body_x[2345] = n_Body_x[2345];
                c_Body_y[2345] = n_Body_y[2345];
                c_Body_x[2346] = n_Body_x[2346];
                c_Body_y[2346] = n_Body_y[2346];
                c_Body_x[2347] = n_Body_x[2347];
                c_Body_y[2347] = n_Body_y[2347];
                c_Body_x[2348] = n_Body_x[2348];
                c_Body_y[2348] = n_Body_y[2348];
                c_Body_x[2349] = n_Body_x[2349];
                c_Body_y[2349] = n_Body_y[2349];
                c_Body_x[2350] = n_Body_x[2350];
                c_Body_y[2350] = n_Body_y[2350];
                c_Body_x[2351] = n_Body_x[2351];
                c_Body_y[2351] = n_Body_y[2351];
                c_Body_x[2352] = n_Body_x[2352];
                c_Body_y[2352] = n_Body_y[2352];
                c_Body_x[2353] = n_Body_x[2353];
                c_Body_y[2353] = n_Body_y[2353];
                c_Body_x[2354] = n_Body_x[2354];
                c_Body_y[2354] = n_Body_y[2354];
                c_Body_x[2355] = n_Body_x[2355];
                c_Body_y[2355] = n_Body_y[2355];
                c_Body_x[2356] = n_Body_x[2356];
                c_Body_y[2356] = n_Body_y[2356];
                c_Body_x[2357] = n_Body_x[2357];
                c_Body_y[2357] = n_Body_y[2357];
                c_Body_x[2358] = n_Body_x[2358];
                c_Body_y[2358] = n_Body_y[2358];
                c_Body_x[2359] = n_Body_x[2359];
                c_Body_y[2359] = n_Body_y[2359];
                c_Body_x[2360] = n_Body_x[2360];
                c_Body_y[2360] = n_Body_y[2360];
                c_Body_x[2361] = n_Body_x[2361];
                c_Body_y[2361] = n_Body_y[2361];
                c_Body_x[2362] = n_Body_x[2362];
                c_Body_y[2362] = n_Body_y[2362];
                c_Body_x[2363] = n_Body_x[2363];
                c_Body_y[2363] = n_Body_y[2363];
                c_Body_x[2364] = n_Body_x[2364];
                c_Body_y[2364] = n_Body_y[2364];
                c_Body_x[2365] = n_Body_x[2365];
                c_Body_y[2365] = n_Body_y[2365];
                c_Body_x[2366] = n_Body_x[2366];
                c_Body_y[2366] = n_Body_y[2366];
                c_Body_x[2367] = n_Body_x[2367];
                c_Body_y[2367] = n_Body_y[2367];
                c_Body_x[2368] = n_Body_x[2368];
                c_Body_y[2368] = n_Body_y[2368];
                c_Body_x[2369] = n_Body_x[2369];
                c_Body_y[2369] = n_Body_y[2369];
                c_Body_x[2370] = n_Body_x[2370];
                c_Body_y[2370] = n_Body_y[2370];
                c_Body_x[2371] = n_Body_x[2371];
                c_Body_y[2371] = n_Body_y[2371];
                c_Body_x[2372] = n_Body_x[2372];
                c_Body_y[2372] = n_Body_y[2372];
                c_Body_x[2373] = n_Body_x[2373];
                c_Body_y[2373] = n_Body_y[2373];
                c_Body_x[2374] = n_Body_x[2374];
                c_Body_y[2374] = n_Body_y[2374];
                c_Body_x[2375] = n_Body_x[2375];
                c_Body_y[2375] = n_Body_y[2375];
                c_Body_x[2376] = n_Body_x[2376];
                c_Body_y[2376] = n_Body_y[2376];
                c_Body_x[2377] = n_Body_x[2377];
                c_Body_y[2377] = n_Body_y[2377];
                c_Body_x[2378] = n_Body_x[2378];
                c_Body_y[2378] = n_Body_y[2378];
                c_Body_x[2379] = n_Body_x[2379];
                c_Body_y[2379] = n_Body_y[2379];
                c_Body_x[2380] = n_Body_x[2380];
                c_Body_y[2380] = n_Body_y[2380];
                c_Body_x[2381] = n_Body_x[2381];
                c_Body_y[2381] = n_Body_y[2381];
                c_Body_x[2382] = n_Body_x[2382];
                c_Body_y[2382] = n_Body_y[2382];
                c_Body_x[2383] = n_Body_x[2383];
                c_Body_y[2383] = n_Body_y[2383];
                c_Body_x[2384] = n_Body_x[2384];
                c_Body_y[2384] = n_Body_y[2384];
                c_Body_x[2385] = n_Body_x[2385];
                c_Body_y[2385] = n_Body_y[2385];
                c_Body_x[2386] = n_Body_x[2386];
                c_Body_y[2386] = n_Body_y[2386];
                c_Body_x[2387] = n_Body_x[2387];
                c_Body_y[2387] = n_Body_y[2387];
                c_Body_x[2388] = n_Body_x[2388];
                c_Body_y[2388] = n_Body_y[2388];
                c_Body_x[2389] = n_Body_x[2389];
                c_Body_y[2389] = n_Body_y[2389];
                c_Body_x[2390] = n_Body_x[2390];
                c_Body_y[2390] = n_Body_y[2390];
                c_Body_x[2391] = n_Body_x[2391];
                c_Body_y[2391] = n_Body_y[2391];
                c_Body_x[2392] = n_Body_x[2392];
                c_Body_y[2392] = n_Body_y[2392];
                c_Body_x[2393] = n_Body_x[2393];
                c_Body_y[2393] = n_Body_y[2393];
                c_Body_x[2394] = n_Body_x[2394];
                c_Body_y[2394] = n_Body_y[2394];
                c_Body_x[2395] = n_Body_x[2395];
                c_Body_y[2395] = n_Body_y[2395];
                c_Body_x[2396] = n_Body_x[2396];
                c_Body_y[2396] = n_Body_y[2396];
                c_Body_x[2397] = n_Body_x[2397];
                c_Body_y[2397] = n_Body_y[2397];
                c_Body_x[2398] = n_Body_x[2398];
                c_Body_y[2398] = n_Body_y[2398];
                c_Body_x[2399] = n_Body_x[2399];
                c_Body_y[2399] = n_Body_y[2399];
                c_Body_x[2400] = n_Body_x[2400];
                c_Body_y[2400] = n_Body_y[2400];
                c_Body_x[2401] = n_Body_x[2401];
                c_Body_y[2401] = n_Body_y[2401];
                c_Body_x[2402] = n_Body_x[2402];
                c_Body_y[2402] = n_Body_y[2402];
                c_Body_x[2403] = n_Body_x[2403];
                c_Body_y[2403] = n_Body_y[2403];
                c_Body_x[2404] = n_Body_x[2404];
                c_Body_y[2404] = n_Body_y[2404];
                c_Body_x[2405] = n_Body_x[2405];
                c_Body_y[2405] = n_Body_y[2405];
                c_Body_x[2406] = n_Body_x[2406];
                c_Body_y[2406] = n_Body_y[2406];
                c_Body_x[2407] = n_Body_x[2407];
                c_Body_y[2407] = n_Body_y[2407];
                c_Body_x[2408] = n_Body_x[2408];
                c_Body_y[2408] = n_Body_y[2408];
                c_Body_x[2409] = n_Body_x[2409];
                c_Body_y[2409] = n_Body_y[2409];
                c_Body_x[2410] = n_Body_x[2410];
                c_Body_y[2410] = n_Body_y[2410];
                c_Body_x[2411] = n_Body_x[2411];
                c_Body_y[2411] = n_Body_y[2411];
                c_Body_x[2412] = n_Body_x[2412];
                c_Body_y[2412] = n_Body_y[2412];
                c_Body_x[2413] = n_Body_x[2413];
                c_Body_y[2413] = n_Body_y[2413];
                c_Body_x[2414] = n_Body_x[2414];
                c_Body_y[2414] = n_Body_y[2414];
                c_Body_x[2415] = n_Body_x[2415];
                c_Body_y[2415] = n_Body_y[2415];
                c_Body_x[2416] = n_Body_x[2416];
                c_Body_y[2416] = n_Body_y[2416];
                c_Body_x[2417] = n_Body_x[2417];
                c_Body_y[2417] = n_Body_y[2417];
                c_Body_x[2418] = n_Body_x[2418];
                c_Body_y[2418] = n_Body_y[2418];
                c_Body_x[2419] = n_Body_x[2419];
                c_Body_y[2419] = n_Body_y[2419];
                c_Body_x[2420] = n_Body_x[2420];
                c_Body_y[2420] = n_Body_y[2420];
                c_Body_x[2421] = n_Body_x[2421];
                c_Body_y[2421] = n_Body_y[2421];
                c_Body_x[2422] = n_Body_x[2422];
                c_Body_y[2422] = n_Body_y[2422];
                c_Body_x[2423] = n_Body_x[2423];
                c_Body_y[2423] = n_Body_y[2423];
                c_Body_x[2424] = n_Body_x[2424];
                c_Body_y[2424] = n_Body_y[2424];
                c_Body_x[2425] = n_Body_x[2425];
                c_Body_y[2425] = n_Body_y[2425];
                c_Body_x[2426] = n_Body_x[2426];
                c_Body_y[2426] = n_Body_y[2426];
                c_Body_x[2427] = n_Body_x[2427];
                c_Body_y[2427] = n_Body_y[2427];
                c_Body_x[2428] = n_Body_x[2428];
                c_Body_y[2428] = n_Body_y[2428];
                c_Body_x[2429] = n_Body_x[2429];
                c_Body_y[2429] = n_Body_y[2429];
                c_Body_x[2430] = n_Body_x[2430];
                c_Body_y[2430] = n_Body_y[2430];
                c_Body_x[2431] = n_Body_x[2431];
                c_Body_y[2431] = n_Body_y[2431];
                c_Body_x[2432] = n_Body_x[2432];
                c_Body_y[2432] = n_Body_y[2432];
                c_Body_x[2433] = n_Body_x[2433];
                c_Body_y[2433] = n_Body_y[2433];
                c_Body_x[2434] = n_Body_x[2434];
                c_Body_y[2434] = n_Body_y[2434];
                c_Body_x[2435] = n_Body_x[2435];
                c_Body_y[2435] = n_Body_y[2435];
                c_Body_x[2436] = n_Body_x[2436];
                c_Body_y[2436] = n_Body_y[2436];
                c_Body_x[2437] = n_Body_x[2437];
                c_Body_y[2437] = n_Body_y[2437];
                c_Body_x[2438] = n_Body_x[2438];
                c_Body_y[2438] = n_Body_y[2438];
                c_Body_x[2439] = n_Body_x[2439];
                c_Body_y[2439] = n_Body_y[2439];
                c_Body_x[2440] = n_Body_x[2440];
                c_Body_y[2440] = n_Body_y[2440];
                c_Body_x[2441] = n_Body_x[2441];
                c_Body_y[2441] = n_Body_y[2441];
                c_Body_x[2442] = n_Body_x[2442];
                c_Body_y[2442] = n_Body_y[2442];
                c_Body_x[2443] = n_Body_x[2443];
                c_Body_y[2443] = n_Body_y[2443];
                c_Body_x[2444] = n_Body_x[2444];
                c_Body_y[2444] = n_Body_y[2444];
                c_Body_x[2445] = n_Body_x[2445];
                c_Body_y[2445] = n_Body_y[2445];
                c_Body_x[2446] = n_Body_x[2446];
                c_Body_y[2446] = n_Body_y[2446];
                c_Body_x[2447] = n_Body_x[2447];
                c_Body_y[2447] = n_Body_y[2447];
                c_Body_x[2448] = n_Body_x[2448];
                c_Body_y[2448] = n_Body_y[2448];
                c_Body_x[2449] = n_Body_x[2449];
                c_Body_y[2449] = n_Body_y[2449];
                c_Body_x[2450] = n_Body_x[2450];
                c_Body_y[2450] = n_Body_y[2450];
                c_Body_x[2451] = n_Body_x[2451];
                c_Body_y[2451] = n_Body_y[2451];
                c_Body_x[2452] = n_Body_x[2452];
                c_Body_y[2452] = n_Body_y[2452];
                c_Body_x[2453] = n_Body_x[2453];
                c_Body_y[2453] = n_Body_y[2453];
                c_Body_x[2454] = n_Body_x[2454];
                c_Body_y[2454] = n_Body_y[2454];
                c_Body_x[2455] = n_Body_x[2455];
                c_Body_y[2455] = n_Body_y[2455];
                c_Body_x[2456] = n_Body_x[2456];
                c_Body_y[2456] = n_Body_y[2456];
                c_Body_x[2457] = n_Body_x[2457];
                c_Body_y[2457] = n_Body_y[2457];
                c_Body_x[2458] = n_Body_x[2458];
                c_Body_y[2458] = n_Body_y[2458];
                c_Body_x[2459] = n_Body_x[2459];
                c_Body_y[2459] = n_Body_y[2459];
                c_Body_x[2460] = n_Body_x[2460];
                c_Body_y[2460] = n_Body_y[2460];
                c_Body_x[2461] = n_Body_x[2461];
                c_Body_y[2461] = n_Body_y[2461];
                c_Body_x[2462] = n_Body_x[2462];
                c_Body_y[2462] = n_Body_y[2462];
                c_Body_x[2463] = n_Body_x[2463];
                c_Body_y[2463] = n_Body_y[2463];
                c_Body_x[2464] = n_Body_x[2464];
                c_Body_y[2464] = n_Body_y[2464];
                c_Body_x[2465] = n_Body_x[2465];
                c_Body_y[2465] = n_Body_y[2465];
                c_Body_x[2466] = n_Body_x[2466];
                c_Body_y[2466] = n_Body_y[2466];
                c_Body_x[2467] = n_Body_x[2467];
                c_Body_y[2467] = n_Body_y[2467];
                c_Body_x[2468] = n_Body_x[2468];
                c_Body_y[2468] = n_Body_y[2468];
                c_Body_x[2469] = n_Body_x[2469];
                c_Body_y[2469] = n_Body_y[2469];
                c_Body_x[2470] = n_Body_x[2470];
                c_Body_y[2470] = n_Body_y[2470];
                c_Body_x[2471] = n_Body_x[2471];
                c_Body_y[2471] = n_Body_y[2471];
                c_Body_x[2472] = n_Body_x[2472];
                c_Body_y[2472] = n_Body_y[2472];
                c_Body_x[2473] = n_Body_x[2473];
                c_Body_y[2473] = n_Body_y[2473];
                c_Body_x[2474] = n_Body_x[2474];
                c_Body_y[2474] = n_Body_y[2474];
                c_Body_x[2475] = n_Body_x[2475];
                c_Body_y[2475] = n_Body_y[2475];
                c_Body_x[2476] = n_Body_x[2476];
                c_Body_y[2476] = n_Body_y[2476];
                c_Body_x[2477] = n_Body_x[2477];
                c_Body_y[2477] = n_Body_y[2477];
                c_Body_x[2478] = n_Body_x[2478];
                c_Body_y[2478] = n_Body_y[2478];
                c_Body_x[2479] = n_Body_x[2479];
                c_Body_y[2479] = n_Body_y[2479];
                c_Body_x[2480] = n_Body_x[2480];
                c_Body_y[2480] = n_Body_y[2480];
                c_Body_x[2481] = n_Body_x[2481];
                c_Body_y[2481] = n_Body_y[2481];
                c_Body_x[2482] = n_Body_x[2482];
                c_Body_y[2482] = n_Body_y[2482];
                c_Body_x[2483] = n_Body_x[2483];
                c_Body_y[2483] = n_Body_y[2483];
                c_Body_x[2484] = n_Body_x[2484];
                c_Body_y[2484] = n_Body_y[2484];
                c_Body_x[2485] = n_Body_x[2485];
                c_Body_y[2485] = n_Body_y[2485];
                c_Body_x[2486] = n_Body_x[2486];
                c_Body_y[2486] = n_Body_y[2486];
                c_Body_x[2487] = n_Body_x[2487];
                c_Body_y[2487] = n_Body_y[2487];
                c_Body_x[2488] = n_Body_x[2488];
                c_Body_y[2488] = n_Body_y[2488];
                c_Body_x[2489] = n_Body_x[2489];
                c_Body_y[2489] = n_Body_y[2489];
                c_Body_x[2490] = n_Body_x[2490];
                c_Body_y[2490] = n_Body_y[2490];
                c_Body_x[2491] = n_Body_x[2491];
                c_Body_y[2491] = n_Body_y[2491];
                c_Body_x[2492] = n_Body_x[2492];
                c_Body_y[2492] = n_Body_y[2492];
                c_Body_x[2493] = n_Body_x[2493];
                c_Body_y[2493] = n_Body_y[2493];
                c_Body_x[2494] = n_Body_x[2494];
                c_Body_y[2494] = n_Body_y[2494];
                c_Body_x[2495] = n_Body_x[2495];
                c_Body_y[2495] = n_Body_y[2495];
                c_Body_x[2496] = n_Body_x[2496];
                c_Body_y[2496] = n_Body_y[2496];
                c_Body_x[2497] = n_Body_x[2497];
                c_Body_y[2497] = n_Body_y[2497];
                c_Body_x[2498] = n_Body_x[2498];
                c_Body_y[2498] = n_Body_y[2498];
                c_Body_x[2499] = n_Body_x[2499];
                c_Body_y[2499] = n_Body_y[2499];
                c_Body_x[2500] = n_Body_x[2500];
                c_Body_y[2500] = n_Body_y[2500];
                c_Body_x[2501] = n_Body_x[2501];
                c_Body_y[2501] = n_Body_y[2501];
                c_Body_x[2502] = n_Body_x[2502];
                c_Body_y[2502] = n_Body_y[2502];
                c_Body_x[2503] = n_Body_x[2503];
                c_Body_y[2503] = n_Body_y[2503];
                c_Body_x[2504] = n_Body_x[2504];
                c_Body_y[2504] = n_Body_y[2504];
                c_Body_x[2505] = n_Body_x[2505];
                c_Body_y[2505] = n_Body_y[2505];
                c_Body_x[2506] = n_Body_x[2506];
                c_Body_y[2506] = n_Body_y[2506];
                c_Body_x[2507] = n_Body_x[2507];
                c_Body_y[2507] = n_Body_y[2507];
                c_Body_x[2508] = n_Body_x[2508];
                c_Body_y[2508] = n_Body_y[2508];
                c_Body_x[2509] = n_Body_x[2509];
                c_Body_y[2509] = n_Body_y[2509];
                c_Body_x[2510] = n_Body_x[2510];
                c_Body_y[2510] = n_Body_y[2510];
                c_Body_x[2511] = n_Body_x[2511];
                c_Body_y[2511] = n_Body_y[2511];
                c_Body_x[2512] = n_Body_x[2512];
                c_Body_y[2512] = n_Body_y[2512];
                c_Body_x[2513] = n_Body_x[2513];
                c_Body_y[2513] = n_Body_y[2513];
                c_Body_x[2514] = n_Body_x[2514];
                c_Body_y[2514] = n_Body_y[2514];
                c_Body_x[2515] = n_Body_x[2515];
                c_Body_y[2515] = n_Body_y[2515];
                c_Body_x[2516] = n_Body_x[2516];
                c_Body_y[2516] = n_Body_y[2516];
                c_Body_x[2517] = n_Body_x[2517];
                c_Body_y[2517] = n_Body_y[2517];
                c_Body_x[2518] = n_Body_x[2518];
                c_Body_y[2518] = n_Body_y[2518];
                c_Body_x[2519] = n_Body_x[2519];
                c_Body_y[2519] = n_Body_y[2519];
                c_Body_x[2520] = n_Body_x[2520];
                c_Body_y[2520] = n_Body_y[2520];
                c_Body_x[2521] = n_Body_x[2521];
                c_Body_y[2521] = n_Body_y[2521];
                c_Body_x[2522] = n_Body_x[2522];
                c_Body_y[2522] = n_Body_y[2522];
                c_Body_x[2523] = n_Body_x[2523];
                c_Body_y[2523] = n_Body_y[2523];
                c_Body_x[2524] = n_Body_x[2524];
                c_Body_y[2524] = n_Body_y[2524];
                c_Body_x[2525] = n_Body_x[2525];
                c_Body_y[2525] = n_Body_y[2525];
                c_Body_x[2526] = n_Body_x[2526];
                c_Body_y[2526] = n_Body_y[2526];
                c_Body_x[2527] = n_Body_x[2527];
                c_Body_y[2527] = n_Body_y[2527];
                c_Body_x[2528] = n_Body_x[2528];
                c_Body_y[2528] = n_Body_y[2528];
                c_Body_x[2529] = n_Body_x[2529];
                c_Body_y[2529] = n_Body_y[2529];
                c_Body_x[2530] = n_Body_x[2530];
                c_Body_y[2530] = n_Body_y[2530];
                c_Body_x[2531] = n_Body_x[2531];
                c_Body_y[2531] = n_Body_y[2531];
                c_Body_x[2532] = n_Body_x[2532];
                c_Body_y[2532] = n_Body_y[2532];
                c_Body_x[2533] = n_Body_x[2533];
                c_Body_y[2533] = n_Body_y[2533];
                c_Body_x[2534] = n_Body_x[2534];
                c_Body_y[2534] = n_Body_y[2534];
                c_Body_x[2535] = n_Body_x[2535];
                c_Body_y[2535] = n_Body_y[2535];
                c_Body_x[2536] = n_Body_x[2536];
                c_Body_y[2536] = n_Body_y[2536];
                c_Body_x[2537] = n_Body_x[2537];
                c_Body_y[2537] = n_Body_y[2537];
                c_Body_x[2538] = n_Body_x[2538];
                c_Body_y[2538] = n_Body_y[2538];
                c_Body_x[2539] = n_Body_x[2539];
                c_Body_y[2539] = n_Body_y[2539];
                c_Body_x[2540] = n_Body_x[2540];
                c_Body_y[2540] = n_Body_y[2540];
                c_Body_x[2541] = n_Body_x[2541];
                c_Body_y[2541] = n_Body_y[2541];
                c_Body_x[2542] = n_Body_x[2542];
                c_Body_y[2542] = n_Body_y[2542];
                c_Body_x[2543] = n_Body_x[2543];
                c_Body_y[2543] = n_Body_y[2543];
                c_Body_x[2544] = n_Body_x[2544];
                c_Body_y[2544] = n_Body_y[2544];
                c_Body_x[2545] = n_Body_x[2545];
                c_Body_y[2545] = n_Body_y[2545];
                c_Body_x[2546] = n_Body_x[2546];
                c_Body_y[2546] = n_Body_y[2546];
                c_Body_x[2547] = n_Body_x[2547];
                c_Body_y[2547] = n_Body_y[2547];
                c_Body_x[2548] = n_Body_x[2548];
                c_Body_y[2548] = n_Body_y[2548];
                c_Body_x[2549] = n_Body_x[2549];
                c_Body_y[2549] = n_Body_y[2549];
                c_Body_x[2550] = n_Body_x[2550];
                c_Body_y[2550] = n_Body_y[2550];
                c_Body_x[2551] = n_Body_x[2551];
                c_Body_y[2551] = n_Body_y[2551];
                c_Body_x[2552] = n_Body_x[2552];
                c_Body_y[2552] = n_Body_y[2552];
                c_Body_x[2553] = n_Body_x[2553];
                c_Body_y[2553] = n_Body_y[2553];
                c_Body_x[2554] = n_Body_x[2554];
                c_Body_y[2554] = n_Body_y[2554];
                c_Body_x[2555] = n_Body_x[2555];
                c_Body_y[2555] = n_Body_y[2555];
                c_Body_x[2556] = n_Body_x[2556];
                c_Body_y[2556] = n_Body_y[2556];
                c_Body_x[2557] = n_Body_x[2557];
                c_Body_y[2557] = n_Body_y[2557];
                c_Body_x[2558] = n_Body_x[2558];
                c_Body_y[2558] = n_Body_y[2558];
                c_Body_x[2559] = n_Body_x[2559];
                c_Body_y[2559] = n_Body_y[2559];
                c_Body_x[2560] = n_Body_x[2560];
                c_Body_y[2560] = n_Body_y[2560];
                c_Body_x[2561] = n_Body_x[2561];
                c_Body_y[2561] = n_Body_y[2561];
                c_Body_x[2562] = n_Body_x[2562];
                c_Body_y[2562] = n_Body_y[2562];
                c_Body_x[2563] = n_Body_x[2563];
                c_Body_y[2563] = n_Body_y[2563];
                c_Body_x[2564] = n_Body_x[2564];
                c_Body_y[2564] = n_Body_y[2564];
                c_Body_x[2565] = n_Body_x[2565];
                c_Body_y[2565] = n_Body_y[2565];
                c_Body_x[2566] = n_Body_x[2566];
                c_Body_y[2566] = n_Body_y[2566];
                c_Body_x[2567] = n_Body_x[2567];
                c_Body_y[2567] = n_Body_y[2567];
                c_Body_x[2568] = n_Body_x[2568];
                c_Body_y[2568] = n_Body_y[2568];
                c_Body_x[2569] = n_Body_x[2569];
                c_Body_y[2569] = n_Body_y[2569];
                c_Body_x[2570] = n_Body_x[2570];
                c_Body_y[2570] = n_Body_y[2570];
                c_Body_x[2571] = n_Body_x[2571];
                c_Body_y[2571] = n_Body_y[2571];
                c_Body_x[2572] = n_Body_x[2572];
                c_Body_y[2572] = n_Body_y[2572];
                c_Body_x[2573] = n_Body_x[2573];
                c_Body_y[2573] = n_Body_y[2573];
                c_Body_x[2574] = n_Body_x[2574];
                c_Body_y[2574] = n_Body_y[2574];
                c_Body_x[2575] = n_Body_x[2575];
                c_Body_y[2575] = n_Body_y[2575];
                c_Body_x[2576] = n_Body_x[2576];
                c_Body_y[2576] = n_Body_y[2576];
                c_Body_x[2577] = n_Body_x[2577];
                c_Body_y[2577] = n_Body_y[2577];
                c_Body_x[2578] = n_Body_x[2578];
                c_Body_y[2578] = n_Body_y[2578];
                c_Body_x[2579] = n_Body_x[2579];
                c_Body_y[2579] = n_Body_y[2579];
                c_Body_x[2580] = n_Body_x[2580];
                c_Body_y[2580] = n_Body_y[2580];
                c_Body_x[2581] = n_Body_x[2581];
                c_Body_y[2581] = n_Body_y[2581];
                c_Body_x[2582] = n_Body_x[2582];
                c_Body_y[2582] = n_Body_y[2582];
                c_Body_x[2583] = n_Body_x[2583];
                c_Body_y[2583] = n_Body_y[2583];
                c_Body_x[2584] = n_Body_x[2584];
                c_Body_y[2584] = n_Body_y[2584];
                c_Body_x[2585] = n_Body_x[2585];
                c_Body_y[2585] = n_Body_y[2585];
                c_Body_x[2586] = n_Body_x[2586];
                c_Body_y[2586] = n_Body_y[2586];
                c_Body_x[2587] = n_Body_x[2587];
                c_Body_y[2587] = n_Body_y[2587];
                c_Body_x[2588] = n_Body_x[2588];
                c_Body_y[2588] = n_Body_y[2588];
                c_Body_x[2589] = n_Body_x[2589];
                c_Body_y[2589] = n_Body_y[2589];
                c_Body_x[2590] = n_Body_x[2590];
                c_Body_y[2590] = n_Body_y[2590];
                c_Body_x[2591] = n_Body_x[2591];
                c_Body_y[2591] = n_Body_y[2591];
                c_Body_x[2592] = n_Body_x[2592];
                c_Body_y[2592] = n_Body_y[2592];
                c_Body_x[2593] = n_Body_x[2593];
                c_Body_y[2593] = n_Body_y[2593];
                c_Body_x[2594] = n_Body_x[2594];
                c_Body_y[2594] = n_Body_y[2594];
                c_Body_x[2595] = n_Body_x[2595];
                c_Body_y[2595] = n_Body_y[2595];
                c_Body_x[2596] = n_Body_x[2596];
                c_Body_y[2596] = n_Body_y[2596];
                c_Body_x[2597] = n_Body_x[2597];
                c_Body_y[2597] = n_Body_y[2597];
                c_Body_x[2598] = n_Body_x[2598];
                c_Body_y[2598] = n_Body_y[2598];
                c_Body_x[2599] = n_Body_x[2599];
                c_Body_y[2599] = n_Body_y[2599];
                c_Body_x[2600] = n_Body_x[2600];
                c_Body_y[2600] = n_Body_y[2600];
                c_Body_x[2601] = n_Body_x[2601];
                c_Body_y[2601] = n_Body_y[2601];
                c_Body_x[2602] = n_Body_x[2602];
                c_Body_y[2602] = n_Body_y[2602];
                c_Body_x[2603] = n_Body_x[2603];
                c_Body_y[2603] = n_Body_y[2603];
                c_Body_x[2604] = n_Body_x[2604];
                c_Body_y[2604] = n_Body_y[2604];
                c_Body_x[2605] = n_Body_x[2605];
                c_Body_y[2605] = n_Body_y[2605];
                c_Body_x[2606] = n_Body_x[2606];
                c_Body_y[2606] = n_Body_y[2606];
                c_Body_x[2607] = n_Body_x[2607];
                c_Body_y[2607] = n_Body_y[2607];
                c_Body_x[2608] = n_Body_x[2608];
                c_Body_y[2608] = n_Body_y[2608];
                c_Body_x[2609] = n_Body_x[2609];
                c_Body_y[2609] = n_Body_y[2609];
                c_Body_x[2610] = n_Body_x[2610];
                c_Body_y[2610] = n_Body_y[2610];
                c_Body_x[2611] = n_Body_x[2611];
                c_Body_y[2611] = n_Body_y[2611];
                c_Body_x[2612] = n_Body_x[2612];
                c_Body_y[2612] = n_Body_y[2612];
                c_Body_x[2613] = n_Body_x[2613];
                c_Body_y[2613] = n_Body_y[2613];
                c_Body_x[2614] = n_Body_x[2614];
                c_Body_y[2614] = n_Body_y[2614];
                c_Body_x[2615] = n_Body_x[2615];
                c_Body_y[2615] = n_Body_y[2615];
                c_Body_x[2616] = n_Body_x[2616];
                c_Body_y[2616] = n_Body_y[2616];
                c_Body_x[2617] = n_Body_x[2617];
                c_Body_y[2617] = n_Body_y[2617];
                c_Body_x[2618] = n_Body_x[2618];
                c_Body_y[2618] = n_Body_y[2618];
                c_Body_x[2619] = n_Body_x[2619];
                c_Body_y[2619] = n_Body_y[2619];
                c_Body_x[2620] = n_Body_x[2620];
                c_Body_y[2620] = n_Body_y[2620];
                c_Body_x[2621] = n_Body_x[2621];
                c_Body_y[2621] = n_Body_y[2621];
                c_Body_x[2622] = n_Body_x[2622];
                c_Body_y[2622] = n_Body_y[2622];
                c_Body_x[2623] = n_Body_x[2623];
                c_Body_y[2623] = n_Body_y[2623];
                c_Body_x[2624] = n_Body_x[2624];
                c_Body_y[2624] = n_Body_y[2624];
                c_Body_x[2625] = n_Body_x[2625];
                c_Body_y[2625] = n_Body_y[2625];
                c_Body_x[2626] = n_Body_x[2626];
                c_Body_y[2626] = n_Body_y[2626];
                c_Body_x[2627] = n_Body_x[2627];
                c_Body_y[2627] = n_Body_y[2627];
                c_Body_x[2628] = n_Body_x[2628];
                c_Body_y[2628] = n_Body_y[2628];
                c_Body_x[2629] = n_Body_x[2629];
                c_Body_y[2629] = n_Body_y[2629];
                c_Body_x[2630] = n_Body_x[2630];
                c_Body_y[2630] = n_Body_y[2630];
                c_Body_x[2631] = n_Body_x[2631];
                c_Body_y[2631] = n_Body_y[2631];
                c_Body_x[2632] = n_Body_x[2632];
                c_Body_y[2632] = n_Body_y[2632];
                c_Body_x[2633] = n_Body_x[2633];
                c_Body_y[2633] = n_Body_y[2633];
                c_Body_x[2634] = n_Body_x[2634];
                c_Body_y[2634] = n_Body_y[2634];
                c_Body_x[2635] = n_Body_x[2635];
                c_Body_y[2635] = n_Body_y[2635];
                c_Body_x[2636] = n_Body_x[2636];
                c_Body_y[2636] = n_Body_y[2636];
                c_Body_x[2637] = n_Body_x[2637];
                c_Body_y[2637] = n_Body_y[2637];
                c_Body_x[2638] = n_Body_x[2638];
                c_Body_y[2638] = n_Body_y[2638];
                c_Body_x[2639] = n_Body_x[2639];
                c_Body_y[2639] = n_Body_y[2639];
                c_Body_x[2640] = n_Body_x[2640];
                c_Body_y[2640] = n_Body_y[2640];
                c_Body_x[2641] = n_Body_x[2641];
                c_Body_y[2641] = n_Body_y[2641];
                c_Body_x[2642] = n_Body_x[2642];
                c_Body_y[2642] = n_Body_y[2642];
                c_Body_x[2643] = n_Body_x[2643];
                c_Body_y[2643] = n_Body_y[2643];
                c_Body_x[2644] = n_Body_x[2644];
                c_Body_y[2644] = n_Body_y[2644];
                c_Body_x[2645] = n_Body_x[2645];
                c_Body_y[2645] = n_Body_y[2645];
                c_Body_x[2646] = n_Body_x[2646];
                c_Body_y[2646] = n_Body_y[2646];
                c_Body_x[2647] = n_Body_x[2647];
                c_Body_y[2647] = n_Body_y[2647];
                c_Body_x[2648] = n_Body_x[2648];
                c_Body_y[2648] = n_Body_y[2648];
                c_Body_x[2649] = n_Body_x[2649];
                c_Body_y[2649] = n_Body_y[2649];
                c_Body_x[2650] = n_Body_x[2650];
                c_Body_y[2650] = n_Body_y[2650];
                c_Body_x[2651] = n_Body_x[2651];
                c_Body_y[2651] = n_Body_y[2651];
                c_Body_x[2652] = n_Body_x[2652];
                c_Body_y[2652] = n_Body_y[2652];
                c_Body_x[2653] = n_Body_x[2653];
                c_Body_y[2653] = n_Body_y[2653];
                c_Body_x[2654] = n_Body_x[2654];
                c_Body_y[2654] = n_Body_y[2654];
                c_Body_x[2655] = n_Body_x[2655];
                c_Body_y[2655] = n_Body_y[2655];
                c_Body_x[2656] = n_Body_x[2656];
                c_Body_y[2656] = n_Body_y[2656];
                c_Body_x[2657] = n_Body_x[2657];
                c_Body_y[2657] = n_Body_y[2657];
                c_Body_x[2658] = n_Body_x[2658];
                c_Body_y[2658] = n_Body_y[2658];
                c_Body_x[2659] = n_Body_x[2659];
                c_Body_y[2659] = n_Body_y[2659];
                c_Body_x[2660] = n_Body_x[2660];
                c_Body_y[2660] = n_Body_y[2660];
                c_Body_x[2661] = n_Body_x[2661];
                c_Body_y[2661] = n_Body_y[2661];
                c_Body_x[2662] = n_Body_x[2662];
                c_Body_y[2662] = n_Body_y[2662];
                c_Body_x[2663] = n_Body_x[2663];
                c_Body_y[2663] = n_Body_y[2663];
                c_Body_x[2664] = n_Body_x[2664];
                c_Body_y[2664] = n_Body_y[2664];
                c_Body_x[2665] = n_Body_x[2665];
                c_Body_y[2665] = n_Body_y[2665];
                c_Body_x[2666] = n_Body_x[2666];
                c_Body_y[2666] = n_Body_y[2666];
                c_Body_x[2667] = n_Body_x[2667];
                c_Body_y[2667] = n_Body_y[2667];
                c_Body_x[2668] = n_Body_x[2668];
                c_Body_y[2668] = n_Body_y[2668];
                c_Body_x[2669] = n_Body_x[2669];
                c_Body_y[2669] = n_Body_y[2669];
                c_Body_x[2670] = n_Body_x[2670];
                c_Body_y[2670] = n_Body_y[2670];
                c_Body_x[2671] = n_Body_x[2671];
                c_Body_y[2671] = n_Body_y[2671];
                c_Body_x[2672] = n_Body_x[2672];
                c_Body_y[2672] = n_Body_y[2672];
                c_Body_x[2673] = n_Body_x[2673];
                c_Body_y[2673] = n_Body_y[2673];
                c_Body_x[2674] = n_Body_x[2674];
                c_Body_y[2674] = n_Body_y[2674];
                c_Body_x[2675] = n_Body_x[2675];
                c_Body_y[2675] = n_Body_y[2675];
                c_Body_x[2676] = n_Body_x[2676];
                c_Body_y[2676] = n_Body_y[2676];
                c_Body_x[2677] = n_Body_x[2677];
                c_Body_y[2677] = n_Body_y[2677];
                c_Body_x[2678] = n_Body_x[2678];
                c_Body_y[2678] = n_Body_y[2678];
                c_Body_x[2679] = n_Body_x[2679];
                c_Body_y[2679] = n_Body_y[2679];
                c_Body_x[2680] = n_Body_x[2680];
                c_Body_y[2680] = n_Body_y[2680];
                c_Body_x[2681] = n_Body_x[2681];
                c_Body_y[2681] = n_Body_y[2681];
                c_Body_x[2682] = n_Body_x[2682];
                c_Body_y[2682] = n_Body_y[2682];
                c_Body_x[2683] = n_Body_x[2683];
                c_Body_y[2683] = n_Body_y[2683];
                c_Body_x[2684] = n_Body_x[2684];
                c_Body_y[2684] = n_Body_y[2684];
                c_Body_x[2685] = n_Body_x[2685];
                c_Body_y[2685] = n_Body_y[2685];
                c_Body_x[2686] = n_Body_x[2686];
                c_Body_y[2686] = n_Body_y[2686];
                c_Body_x[2687] = n_Body_x[2687];
                c_Body_y[2687] = n_Body_y[2687];
                c_Body_x[2688] = n_Body_x[2688];
                c_Body_y[2688] = n_Body_y[2688];
                c_Body_x[2689] = n_Body_x[2689];
                c_Body_y[2689] = n_Body_y[2689];
                c_Body_x[2690] = n_Body_x[2690];
                c_Body_y[2690] = n_Body_y[2690];
                c_Body_x[2691] = n_Body_x[2691];
                c_Body_y[2691] = n_Body_y[2691];
                c_Body_x[2692] = n_Body_x[2692];
                c_Body_y[2692] = n_Body_y[2692];
                c_Body_x[2693] = n_Body_x[2693];
                c_Body_y[2693] = n_Body_y[2693];
                c_Body_x[2694] = n_Body_x[2694];
                c_Body_y[2694] = n_Body_y[2694];
                c_Body_x[2695] = n_Body_x[2695];
                c_Body_y[2695] = n_Body_y[2695];
                c_Body_x[2696] = n_Body_x[2696];
                c_Body_y[2696] = n_Body_y[2696];
                c_Body_x[2697] = n_Body_x[2697];
                c_Body_y[2697] = n_Body_y[2697];
                c_Body_x[2698] = n_Body_x[2698];
                c_Body_y[2698] = n_Body_y[2698];
                c_Body_x[2699] = n_Body_x[2699];
                c_Body_y[2699] = n_Body_y[2699];
                c_Body_x[2700] = n_Body_x[2700];
                c_Body_y[2700] = n_Body_y[2700];
                c_Body_x[2701] = n_Body_x[2701];
                c_Body_y[2701] = n_Body_y[2701];
                c_Body_x[2702] = n_Body_x[2702];
                c_Body_y[2702] = n_Body_y[2702];
                c_Body_x[2703] = n_Body_x[2703];
                c_Body_y[2703] = n_Body_y[2703];
                c_Body_x[2704] = n_Body_x[2704];
                c_Body_y[2704] = n_Body_y[2704];
                c_Body_x[2705] = n_Body_x[2705];
                c_Body_y[2705] = n_Body_y[2705];
                c_Body_x[2706] = n_Body_x[2706];
                c_Body_y[2706] = n_Body_y[2706];
                c_Body_x[2707] = n_Body_x[2707];
                c_Body_y[2707] = n_Body_y[2707];
                c_Body_x[2708] = n_Body_x[2708];
                c_Body_y[2708] = n_Body_y[2708];
                c_Body_x[2709] = n_Body_x[2709];
                c_Body_y[2709] = n_Body_y[2709];
                c_Body_x[2710] = n_Body_x[2710];
                c_Body_y[2710] = n_Body_y[2710];
                c_Body_x[2711] = n_Body_x[2711];
                c_Body_y[2711] = n_Body_y[2711];
                c_Body_x[2712] = n_Body_x[2712];
                c_Body_y[2712] = n_Body_y[2712];
                c_Body_x[2713] = n_Body_x[2713];
                c_Body_y[2713] = n_Body_y[2713];
                c_Body_x[2714] = n_Body_x[2714];
                c_Body_y[2714] = n_Body_y[2714];
                c_Body_x[2715] = n_Body_x[2715];
                c_Body_y[2715] = n_Body_y[2715];
                c_Body_x[2716] = n_Body_x[2716];
                c_Body_y[2716] = n_Body_y[2716];
                c_Body_x[2717] = n_Body_x[2717];
                c_Body_y[2717] = n_Body_y[2717];
                c_Body_x[2718] = n_Body_x[2718];
                c_Body_y[2718] = n_Body_y[2718];
                c_Body_x[2719] = n_Body_x[2719];
                c_Body_y[2719] = n_Body_y[2719];
                c_Body_x[2720] = n_Body_x[2720];
                c_Body_y[2720] = n_Body_y[2720];
                c_Body_x[2721] = n_Body_x[2721];
                c_Body_y[2721] = n_Body_y[2721];
                c_Body_x[2722] = n_Body_x[2722];
                c_Body_y[2722] = n_Body_y[2722];
                c_Body_x[2723] = n_Body_x[2723];
                c_Body_y[2723] = n_Body_y[2723];
                c_Body_x[2724] = n_Body_x[2724];
                c_Body_y[2724] = n_Body_y[2724];
                c_Body_x[2725] = n_Body_x[2725];
                c_Body_y[2725] = n_Body_y[2725];
                c_Body_x[2726] = n_Body_x[2726];
                c_Body_y[2726] = n_Body_y[2726];
                c_Body_x[2727] = n_Body_x[2727];
                c_Body_y[2727] = n_Body_y[2727];
                c_Body_x[2728] = n_Body_x[2728];
                c_Body_y[2728] = n_Body_y[2728];
                c_Body_x[2729] = n_Body_x[2729];
                c_Body_y[2729] = n_Body_y[2729];
                c_Body_x[2730] = n_Body_x[2730];
                c_Body_y[2730] = n_Body_y[2730];
                c_Body_x[2731] = n_Body_x[2731];
                c_Body_y[2731] = n_Body_y[2731];
                c_Body_x[2732] = n_Body_x[2732];
                c_Body_y[2732] = n_Body_y[2732];
                c_Body_x[2733] = n_Body_x[2733];
                c_Body_y[2733] = n_Body_y[2733];
                c_Body_x[2734] = n_Body_x[2734];
                c_Body_y[2734] = n_Body_y[2734];
                c_Body_x[2735] = n_Body_x[2735];
                c_Body_y[2735] = n_Body_y[2735];
                c_Body_x[2736] = n_Body_x[2736];
                c_Body_y[2736] = n_Body_y[2736];
                c_Body_x[2737] = n_Body_x[2737];
                c_Body_y[2737] = n_Body_y[2737];
                c_Body_x[2738] = n_Body_x[2738];
                c_Body_y[2738] = n_Body_y[2738];
                c_Body_x[2739] = n_Body_x[2739];
                c_Body_y[2739] = n_Body_y[2739];
                c_Body_x[2740] = n_Body_x[2740];
                c_Body_y[2740] = n_Body_y[2740];
                c_Body_x[2741] = n_Body_x[2741];
                c_Body_y[2741] = n_Body_y[2741];
                c_Body_x[2742] = n_Body_x[2742];
                c_Body_y[2742] = n_Body_y[2742];
                c_Body_x[2743] = n_Body_x[2743];
                c_Body_y[2743] = n_Body_y[2743];
                c_Body_x[2744] = n_Body_x[2744];
                c_Body_y[2744] = n_Body_y[2744];
                c_Body_x[2745] = n_Body_x[2745];
                c_Body_y[2745] = n_Body_y[2745];
                c_Body_x[2746] = n_Body_x[2746];
                c_Body_y[2746] = n_Body_y[2746];
                c_Body_x[2747] = n_Body_x[2747];
                c_Body_y[2747] = n_Body_y[2747];
                c_Body_x[2748] = n_Body_x[2748];
                c_Body_y[2748] = n_Body_y[2748];
                c_Body_x[2749] = n_Body_x[2749];
                c_Body_y[2749] = n_Body_y[2749];
                c_Body_x[2750] = n_Body_x[2750];
                c_Body_y[2750] = n_Body_y[2750];
                c_Body_x[2751] = n_Body_x[2751];
                c_Body_y[2751] = n_Body_y[2751];
                c_Body_x[2752] = n_Body_x[2752];
                c_Body_y[2752] = n_Body_y[2752];
                c_Body_x[2753] = n_Body_x[2753];
                c_Body_y[2753] = n_Body_y[2753];
                c_Body_x[2754] = n_Body_x[2754];
                c_Body_y[2754] = n_Body_y[2754];
                c_Body_x[2755] = n_Body_x[2755];
                c_Body_y[2755] = n_Body_y[2755];
                c_Body_x[2756] = n_Body_x[2756];
                c_Body_y[2756] = n_Body_y[2756];
                c_Body_x[2757] = n_Body_x[2757];
                c_Body_y[2757] = n_Body_y[2757];
                c_Body_x[2758] = n_Body_x[2758];
                c_Body_y[2758] = n_Body_y[2758];
                c_Body_x[2759] = n_Body_x[2759];
                c_Body_y[2759] = n_Body_y[2759];
                c_Body_x[2760] = n_Body_x[2760];
                c_Body_y[2760] = n_Body_y[2760];
                c_Body_x[2761] = n_Body_x[2761];
                c_Body_y[2761] = n_Body_y[2761];
                c_Body_x[2762] = n_Body_x[2762];
                c_Body_y[2762] = n_Body_y[2762];
                c_Body_x[2763] = n_Body_x[2763];
                c_Body_y[2763] = n_Body_y[2763];
                c_Body_x[2764] = n_Body_x[2764];
                c_Body_y[2764] = n_Body_y[2764];
                c_Body_x[2765] = n_Body_x[2765];
                c_Body_y[2765] = n_Body_y[2765];
                c_Body_x[2766] = n_Body_x[2766];
                c_Body_y[2766] = n_Body_y[2766];
                c_Body_x[2767] = n_Body_x[2767];
                c_Body_y[2767] = n_Body_y[2767];
                c_Body_x[2768] = n_Body_x[2768];
                c_Body_y[2768] = n_Body_y[2768];
                c_Body_x[2769] = n_Body_x[2769];
                c_Body_y[2769] = n_Body_y[2769];
                c_Body_x[2770] = n_Body_x[2770];
                c_Body_y[2770] = n_Body_y[2770];
                c_Body_x[2771] = n_Body_x[2771];
                c_Body_y[2771] = n_Body_y[2771];
                c_Body_x[2772] = n_Body_x[2772];
                c_Body_y[2772] = n_Body_y[2772];
                c_Body_x[2773] = n_Body_x[2773];
                c_Body_y[2773] = n_Body_y[2773];
                c_Body_x[2774] = n_Body_x[2774];
                c_Body_y[2774] = n_Body_y[2774];
                c_Body_x[2775] = n_Body_x[2775];
                c_Body_y[2775] = n_Body_y[2775];
                c_Body_x[2776] = n_Body_x[2776];
                c_Body_y[2776] = n_Body_y[2776];
                c_Body_x[2777] = n_Body_x[2777];
                c_Body_y[2777] = n_Body_y[2777];
                c_Body_x[2778] = n_Body_x[2778];
                c_Body_y[2778] = n_Body_y[2778];
                c_Body_x[2779] = n_Body_x[2779];
                c_Body_y[2779] = n_Body_y[2779];
                c_Body_x[2780] = n_Body_x[2780];
                c_Body_y[2780] = n_Body_y[2780];
                c_Body_x[2781] = n_Body_x[2781];
                c_Body_y[2781] = n_Body_y[2781];
                c_Body_x[2782] = n_Body_x[2782];
                c_Body_y[2782] = n_Body_y[2782];
                c_Body_x[2783] = n_Body_x[2783];
                c_Body_y[2783] = n_Body_y[2783];
                c_Body_x[2784] = n_Body_x[2784];
                c_Body_y[2784] = n_Body_y[2784];
                c_Body_x[2785] = n_Body_x[2785];
                c_Body_y[2785] = n_Body_y[2785];
                c_Body_x[2786] = n_Body_x[2786];
                c_Body_y[2786] = n_Body_y[2786];
                c_Body_x[2787] = n_Body_x[2787];
                c_Body_y[2787] = n_Body_y[2787];
                c_Body_x[2788] = n_Body_x[2788];
                c_Body_y[2788] = n_Body_y[2788];
                c_Body_x[2789] = n_Body_x[2789];
                c_Body_y[2789] = n_Body_y[2789];
                c_Body_x[2790] = n_Body_x[2790];
                c_Body_y[2790] = n_Body_y[2790];
                c_Body_x[2791] = n_Body_x[2791];
                c_Body_y[2791] = n_Body_y[2791];
                c_Body_x[2792] = n_Body_x[2792];
                c_Body_y[2792] = n_Body_y[2792];
                c_Body_x[2793] = n_Body_x[2793];
                c_Body_y[2793] = n_Body_y[2793];
                c_Body_x[2794] = n_Body_x[2794];
                c_Body_y[2794] = n_Body_y[2794];
                c_Body_x[2795] = n_Body_x[2795];
                c_Body_y[2795] = n_Body_y[2795];
                c_Body_x[2796] = n_Body_x[2796];
                c_Body_y[2796] = n_Body_y[2796];
                c_Body_x[2797] = n_Body_x[2797];
                c_Body_y[2797] = n_Body_y[2797];
                c_Body_x[2798] = n_Body_x[2798];
                c_Body_y[2798] = n_Body_y[2798];
                c_Body_x[2799] = n_Body_x[2799];
                c_Body_y[2799] = n_Body_y[2799];
                c_Body_x[2800] = n_Body_x[2800];
                c_Body_y[2800] = n_Body_y[2800];
                c_Body_x[2801] = n_Body_x[2801];
                c_Body_y[2801] = n_Body_y[2801];
                c_Body_x[2802] = n_Body_x[2802];
                c_Body_y[2802] = n_Body_y[2802];
                c_Body_x[2803] = n_Body_x[2803];
                c_Body_y[2803] = n_Body_y[2803];
                c_Body_x[2804] = n_Body_x[2804];
                c_Body_y[2804] = n_Body_y[2804];
                c_Body_x[2805] = n_Body_x[2805];
                c_Body_y[2805] = n_Body_y[2805];
                c_Body_x[2806] = n_Body_x[2806];
                c_Body_y[2806] = n_Body_y[2806];
                c_Body_x[2807] = n_Body_x[2807];
                c_Body_y[2807] = n_Body_y[2807];
                c_Body_x[2808] = n_Body_x[2808];
                c_Body_y[2808] = n_Body_y[2808];
                c_Body_x[2809] = n_Body_x[2809];
                c_Body_y[2809] = n_Body_y[2809];
                c_Body_x[2810] = n_Body_x[2810];
                c_Body_y[2810] = n_Body_y[2810];
                c_Body_x[2811] = n_Body_x[2811];
                c_Body_y[2811] = n_Body_y[2811];
                c_Body_x[2812] = n_Body_x[2812];
                c_Body_y[2812] = n_Body_y[2812];
                c_Body_x[2813] = n_Body_x[2813];
                c_Body_y[2813] = n_Body_y[2813];
                c_Body_x[2814] = n_Body_x[2814];
                c_Body_y[2814] = n_Body_y[2814];
                c_Body_x[2815] = n_Body_x[2815];
                c_Body_y[2815] = n_Body_y[2815];
                c_Body_x[2816] = n_Body_x[2816];
                c_Body_y[2816] = n_Body_y[2816];
                c_Body_x[2817] = n_Body_x[2817];
                c_Body_y[2817] = n_Body_y[2817];
                c_Body_x[2818] = n_Body_x[2818];
                c_Body_y[2818] = n_Body_y[2818];
                c_Body_x[2819] = n_Body_x[2819];
                c_Body_y[2819] = n_Body_y[2819];
                c_Body_x[2820] = n_Body_x[2820];
                c_Body_y[2820] = n_Body_y[2820];
                c_Body_x[2821] = n_Body_x[2821];
                c_Body_y[2821] = n_Body_y[2821];
                c_Body_x[2822] = n_Body_x[2822];
                c_Body_y[2822] = n_Body_y[2822];
                c_Body_x[2823] = n_Body_x[2823];
                c_Body_y[2823] = n_Body_y[2823];
                c_Body_x[2824] = n_Body_x[2824];
                c_Body_y[2824] = n_Body_y[2824];
                c_Body_x[2825] = n_Body_x[2825];
                c_Body_y[2825] = n_Body_y[2825];
                c_Body_x[2826] = n_Body_x[2826];
                c_Body_y[2826] = n_Body_y[2826];
                c_Body_x[2827] = n_Body_x[2827];
                c_Body_y[2827] = n_Body_y[2827];
                c_Body_x[2828] = n_Body_x[2828];
                c_Body_y[2828] = n_Body_y[2828];
                c_Body_x[2829] = n_Body_x[2829];
                c_Body_y[2829] = n_Body_y[2829];
                c_Body_x[2830] = n_Body_x[2830];
                c_Body_y[2830] = n_Body_y[2830];
                c_Body_x[2831] = n_Body_x[2831];
                c_Body_y[2831] = n_Body_y[2831];
                c_Body_x[2832] = n_Body_x[2832];
                c_Body_y[2832] = n_Body_y[2832];
                c_Body_x[2833] = n_Body_x[2833];
                c_Body_y[2833] = n_Body_y[2833];
                c_Body_x[2834] = n_Body_x[2834];
                c_Body_y[2834] = n_Body_y[2834];
                c_Body_x[2835] = n_Body_x[2835];
                c_Body_y[2835] = n_Body_y[2835];
                c_Body_x[2836] = n_Body_x[2836];
                c_Body_y[2836] = n_Body_y[2836];
                c_Body_x[2837] = n_Body_x[2837];
                c_Body_y[2837] = n_Body_y[2837];
                c_Body_x[2838] = n_Body_x[2838];
                c_Body_y[2838] = n_Body_y[2838];
                c_Body_x[2839] = n_Body_x[2839];
                c_Body_y[2839] = n_Body_y[2839];
                c_Body_x[2840] = n_Body_x[2840];
                c_Body_y[2840] = n_Body_y[2840];
                c_Body_x[2841] = n_Body_x[2841];
                c_Body_y[2841] = n_Body_y[2841];
                c_Body_x[2842] = n_Body_x[2842];
                c_Body_y[2842] = n_Body_y[2842];
                c_Body_x[2843] = n_Body_x[2843];
                c_Body_y[2843] = n_Body_y[2843];
                c_Body_x[2844] = n_Body_x[2844];
                c_Body_y[2844] = n_Body_y[2844];
                c_Body_x[2845] = n_Body_x[2845];
                c_Body_y[2845] = n_Body_y[2845];
                c_Body_x[2846] = n_Body_x[2846];
                c_Body_y[2846] = n_Body_y[2846];
                c_Body_x[2847] = n_Body_x[2847];
                c_Body_y[2847] = n_Body_y[2847];
                c_Body_x[2848] = n_Body_x[2848];
                c_Body_y[2848] = n_Body_y[2848];
                c_Body_x[2849] = n_Body_x[2849];
                c_Body_y[2849] = n_Body_y[2849];
                c_Body_x[2850] = n_Body_x[2850];
                c_Body_y[2850] = n_Body_y[2850];
                c_Body_x[2851] = n_Body_x[2851];
                c_Body_y[2851] = n_Body_y[2851];
                c_Body_x[2852] = n_Body_x[2852];
                c_Body_y[2852] = n_Body_y[2852];
                c_Body_x[2853] = n_Body_x[2853];
                c_Body_y[2853] = n_Body_y[2853];
                c_Body_x[2854] = n_Body_x[2854];
                c_Body_y[2854] = n_Body_y[2854];
                c_Body_x[2855] = n_Body_x[2855];
                c_Body_y[2855] = n_Body_y[2855];
                c_Body_x[2856] = n_Body_x[2856];
                c_Body_y[2856] = n_Body_y[2856];
                c_Body_x[2857] = n_Body_x[2857];
                c_Body_y[2857] = n_Body_y[2857];
                c_Body_x[2858] = n_Body_x[2858];
                c_Body_y[2858] = n_Body_y[2858];
                c_Body_x[2859] = n_Body_x[2859];
                c_Body_y[2859] = n_Body_y[2859];
                c_Body_x[2860] = n_Body_x[2860];
                c_Body_y[2860] = n_Body_y[2860];
                c_Body_x[2861] = n_Body_x[2861];
                c_Body_y[2861] = n_Body_y[2861];
                c_Body_x[2862] = n_Body_x[2862];
                c_Body_y[2862] = n_Body_y[2862];
                c_Body_x[2863] = n_Body_x[2863];
                c_Body_y[2863] = n_Body_y[2863];
                c_Body_x[2864] = n_Body_x[2864];
                c_Body_y[2864] = n_Body_y[2864];
                c_Body_x[2865] = n_Body_x[2865];
                c_Body_y[2865] = n_Body_y[2865];
                c_Body_x[2866] = n_Body_x[2866];
                c_Body_y[2866] = n_Body_y[2866];
                c_Body_x[2867] = n_Body_x[2867];
                c_Body_y[2867] = n_Body_y[2867];
                c_Body_x[2868] = n_Body_x[2868];
                c_Body_y[2868] = n_Body_y[2868];
                c_Body_x[2869] = n_Body_x[2869];
                c_Body_y[2869] = n_Body_y[2869];
                c_Body_x[2870] = n_Body_x[2870];
                c_Body_y[2870] = n_Body_y[2870];
                c_Body_x[2871] = n_Body_x[2871];
                c_Body_y[2871] = n_Body_y[2871];
                c_Body_x[2872] = n_Body_x[2872];
                c_Body_y[2872] = n_Body_y[2872];
                c_Body_x[2873] = n_Body_x[2873];
                c_Body_y[2873] = n_Body_y[2873];
                c_Body_x[2874] = n_Body_x[2874];
                c_Body_y[2874] = n_Body_y[2874];
                c_Body_x[2875] = n_Body_x[2875];
                c_Body_y[2875] = n_Body_y[2875];
                c_Body_x[2876] = n_Body_x[2876];
                c_Body_y[2876] = n_Body_y[2876];
                c_Body_x[2877] = n_Body_x[2877];
                c_Body_y[2877] = n_Body_y[2877];
                c_Body_x[2878] = n_Body_x[2878];
                c_Body_y[2878] = n_Body_y[2878];
                c_Body_x[2879] = n_Body_x[2879];
                c_Body_y[2879] = n_Body_y[2879];
                c_Body_x[2880] = n_Body_x[2880];
                c_Body_y[2880] = n_Body_y[2880];
                c_Body_x[2881] = n_Body_x[2881];
                c_Body_y[2881] = n_Body_y[2881];
                c_Body_x[2882] = n_Body_x[2882];
                c_Body_y[2882] = n_Body_y[2882];
                c_Body_x[2883] = n_Body_x[2883];
                c_Body_y[2883] = n_Body_y[2883];
                c_Body_x[2884] = n_Body_x[2884];
                c_Body_y[2884] = n_Body_y[2884];
                c_Body_x[2885] = n_Body_x[2885];
                c_Body_y[2885] = n_Body_y[2885];
                c_Body_x[2886] = n_Body_x[2886];
                c_Body_y[2886] = n_Body_y[2886];
                c_Body_x[2887] = n_Body_x[2887];
                c_Body_y[2887] = n_Body_y[2887];
                c_Body_x[2888] = n_Body_x[2888];
                c_Body_y[2888] = n_Body_y[2888];
                c_Body_x[2889] = n_Body_x[2889];
                c_Body_y[2889] = n_Body_y[2889];
                c_Body_x[2890] = n_Body_x[2890];
                c_Body_y[2890] = n_Body_y[2890];
                c_Body_x[2891] = n_Body_x[2891];
                c_Body_y[2891] = n_Body_y[2891];
                c_Body_x[2892] = n_Body_x[2892];
                c_Body_y[2892] = n_Body_y[2892];
                c_Body_x[2893] = n_Body_x[2893];
                c_Body_y[2893] = n_Body_y[2893];
                c_Body_x[2894] = n_Body_x[2894];
                c_Body_y[2894] = n_Body_y[2894];
                c_Body_x[2895] = n_Body_x[2895];
                c_Body_y[2895] = n_Body_y[2895];
                c_Body_x[2896] = n_Body_x[2896];
                c_Body_y[2896] = n_Body_y[2896];
                c_Body_x[2897] = n_Body_x[2897];
                c_Body_y[2897] = n_Body_y[2897];
                c_Body_x[2898] = n_Body_x[2898];
                c_Body_y[2898] = n_Body_y[2898];
                c_Body_x[2899] = n_Body_x[2899];
                c_Body_y[2899] = n_Body_y[2899];
                c_Body_x[2900] = n_Body_x[2900];
                c_Body_y[2900] = n_Body_y[2900];
                c_Body_x[2901] = n_Body_x[2901];
                c_Body_y[2901] = n_Body_y[2901];
                c_Body_x[2902] = n_Body_x[2902];
                c_Body_y[2902] = n_Body_y[2902];
                c_Body_x[2903] = n_Body_x[2903];
                c_Body_y[2903] = n_Body_y[2903];
                c_Body_x[2904] = n_Body_x[2904];
                c_Body_y[2904] = n_Body_y[2904];
                c_Body_x[2905] = n_Body_x[2905];
                c_Body_y[2905] = n_Body_y[2905];
                c_Body_x[2906] = n_Body_x[2906];
                c_Body_y[2906] = n_Body_y[2906];
                c_Body_x[2907] = n_Body_x[2907];
                c_Body_y[2907] = n_Body_y[2907];
                c_Body_x[2908] = n_Body_x[2908];
                c_Body_y[2908] = n_Body_y[2908];
                c_Body_x[2909] = n_Body_x[2909];
                c_Body_y[2909] = n_Body_y[2909];
                c_Body_x[2910] = n_Body_x[2910];
                c_Body_y[2910] = n_Body_y[2910];
                c_Body_x[2911] = n_Body_x[2911];
                c_Body_y[2911] = n_Body_y[2911];
                c_Body_x[2912] = n_Body_x[2912];
                c_Body_y[2912] = n_Body_y[2912];
                c_Body_x[2913] = n_Body_x[2913];
                c_Body_y[2913] = n_Body_y[2913];
                c_Body_x[2914] = n_Body_x[2914];
                c_Body_y[2914] = n_Body_y[2914];
                c_Body_x[2915] = n_Body_x[2915];
                c_Body_y[2915] = n_Body_y[2915];
                c_Body_x[2916] = n_Body_x[2916];
                c_Body_y[2916] = n_Body_y[2916];
                c_Body_x[2917] = n_Body_x[2917];
                c_Body_y[2917] = n_Body_y[2917];
                c_Body_x[2918] = n_Body_x[2918];
                c_Body_y[2918] = n_Body_y[2918];
                c_Body_x[2919] = n_Body_x[2919];
                c_Body_y[2919] = n_Body_y[2919];
                c_Body_x[2920] = n_Body_x[2920];
                c_Body_y[2920] = n_Body_y[2920];
                c_Body_x[2921] = n_Body_x[2921];
                c_Body_y[2921] = n_Body_y[2921];
                c_Body_x[2922] = n_Body_x[2922];
                c_Body_y[2922] = n_Body_y[2922];
                c_Body_x[2923] = n_Body_x[2923];
                c_Body_y[2923] = n_Body_y[2923];
                c_Body_x[2924] = n_Body_x[2924];
                c_Body_y[2924] = n_Body_y[2924];
                c_Body_x[2925] = n_Body_x[2925];
                c_Body_y[2925] = n_Body_y[2925];
                c_Body_x[2926] = n_Body_x[2926];
                c_Body_y[2926] = n_Body_y[2926];
                c_Body_x[2927] = n_Body_x[2927];
                c_Body_y[2927] = n_Body_y[2927];
                c_Body_x[2928] = n_Body_x[2928];
                c_Body_y[2928] = n_Body_y[2928];
                c_Body_x[2929] = n_Body_x[2929];
                c_Body_y[2929] = n_Body_y[2929];
                c_Body_x[2930] = n_Body_x[2930];
                c_Body_y[2930] = n_Body_y[2930];
                c_Body_x[2931] = n_Body_x[2931];
                c_Body_y[2931] = n_Body_y[2931];
                c_Body_x[2932] = n_Body_x[2932];
                c_Body_y[2932] = n_Body_y[2932];
                c_Body_x[2933] = n_Body_x[2933];
                c_Body_y[2933] = n_Body_y[2933];
                c_Body_x[2934] = n_Body_x[2934];
                c_Body_y[2934] = n_Body_y[2934];
                c_Body_x[2935] = n_Body_x[2935];
                c_Body_y[2935] = n_Body_y[2935];
                c_Body_x[2936] = n_Body_x[2936];
                c_Body_y[2936] = n_Body_y[2936];
                c_Body_x[2937] = n_Body_x[2937];
                c_Body_y[2937] = n_Body_y[2937];
                c_Body_x[2938] = n_Body_x[2938];
                c_Body_y[2938] = n_Body_y[2938];
                c_Body_x[2939] = n_Body_x[2939];
                c_Body_y[2939] = n_Body_y[2939];
                c_Body_x[2940] = n_Body_x[2940];
                c_Body_y[2940] = n_Body_y[2940];
                c_Body_x[2941] = n_Body_x[2941];
                c_Body_y[2941] = n_Body_y[2941];
                c_Body_x[2942] = n_Body_x[2942];
                c_Body_y[2942] = n_Body_y[2942];
                c_Body_x[2943] = n_Body_x[2943];
                c_Body_y[2943] = n_Body_y[2943];
                c_Body_x[2944] = n_Body_x[2944];
                c_Body_y[2944] = n_Body_y[2944];
                c_Body_x[2945] = n_Body_x[2945];
                c_Body_y[2945] = n_Body_y[2945];
                c_Body_x[2946] = n_Body_x[2946];
                c_Body_y[2946] = n_Body_y[2946];
                c_Body_x[2947] = n_Body_x[2947];
                c_Body_y[2947] = n_Body_y[2947];
                c_Body_x[2948] = n_Body_x[2948];
                c_Body_y[2948] = n_Body_y[2948];
                c_Body_x[2949] = n_Body_x[2949];
                c_Body_y[2949] = n_Body_y[2949];
                c_Body_x[2950] = n_Body_x[2950];
                c_Body_y[2950] = n_Body_y[2950];
                c_Body_x[2951] = n_Body_x[2951];
                c_Body_y[2951] = n_Body_y[2951];
                c_Body_x[2952] = n_Body_x[2952];
                c_Body_y[2952] = n_Body_y[2952];
                c_Body_x[2953] = n_Body_x[2953];
                c_Body_y[2953] = n_Body_y[2953];
                c_Body_x[2954] = n_Body_x[2954];
                c_Body_y[2954] = n_Body_y[2954];
                c_Body_x[2955] = n_Body_x[2955];
                c_Body_y[2955] = n_Body_y[2955];
                c_Body_x[2956] = n_Body_x[2956];
                c_Body_y[2956] = n_Body_y[2956];
                c_Body_x[2957] = n_Body_x[2957];
                c_Body_y[2957] = n_Body_y[2957];
                c_Body_x[2958] = n_Body_x[2958];
                c_Body_y[2958] = n_Body_y[2958];
                c_Body_x[2959] = n_Body_x[2959];
                c_Body_y[2959] = n_Body_y[2959];
                c_Body_x[2960] = n_Body_x[2960];
                c_Body_y[2960] = n_Body_y[2960];
                c_Body_x[2961] = n_Body_x[2961];
                c_Body_y[2961] = n_Body_y[2961];
                c_Body_x[2962] = n_Body_x[2962];
                c_Body_y[2962] = n_Body_y[2962];
                c_Body_x[2963] = n_Body_x[2963];
                c_Body_y[2963] = n_Body_y[2963];
                c_Body_x[2964] = n_Body_x[2964];
                c_Body_y[2964] = n_Body_y[2964];
                c_Body_x[2965] = n_Body_x[2965];
                c_Body_y[2965] = n_Body_y[2965];
                c_Body_x[2966] = n_Body_x[2966];
                c_Body_y[2966] = n_Body_y[2966];
                c_Body_x[2967] = n_Body_x[2967];
                c_Body_y[2967] = n_Body_y[2967];
                c_Body_x[2968] = n_Body_x[2968];
                c_Body_y[2968] = n_Body_y[2968];
                c_Body_x[2969] = n_Body_x[2969];
                c_Body_y[2969] = n_Body_y[2969];
                c_Body_x[2970] = n_Body_x[2970];
                c_Body_y[2970] = n_Body_y[2970];
                c_Body_x[2971] = n_Body_x[2971];
                c_Body_y[2971] = n_Body_y[2971];
                c_Body_x[2972] = n_Body_x[2972];
                c_Body_y[2972] = n_Body_y[2972];
                c_Body_x[2973] = n_Body_x[2973];
                c_Body_y[2973] = n_Body_y[2973];
                c_Body_x[2974] = n_Body_x[2974];
                c_Body_y[2974] = n_Body_y[2974];
                c_Body_x[2975] = n_Body_x[2975];
                c_Body_y[2975] = n_Body_y[2975];
                c_Body_x[2976] = n_Body_x[2976];
                c_Body_y[2976] = n_Body_y[2976];
                c_Body_x[2977] = n_Body_x[2977];
                c_Body_y[2977] = n_Body_y[2977];
                c_Body_x[2978] = n_Body_x[2978];
                c_Body_y[2978] = n_Body_y[2978];
                c_Body_x[2979] = n_Body_x[2979];
                c_Body_y[2979] = n_Body_y[2979];
                c_Body_x[2980] = n_Body_x[2980];
                c_Body_y[2980] = n_Body_y[2980];
                c_Body_x[2981] = n_Body_x[2981];
                c_Body_y[2981] = n_Body_y[2981];
                c_Body_x[2982] = n_Body_x[2982];
                c_Body_y[2982] = n_Body_y[2982];
                c_Body_x[2983] = n_Body_x[2983];
                c_Body_y[2983] = n_Body_y[2983];
                c_Body_x[2984] = n_Body_x[2984];
                c_Body_y[2984] = n_Body_y[2984];
                c_Body_x[2985] = n_Body_x[2985];
                c_Body_y[2985] = n_Body_y[2985];
                c_Body_x[2986] = n_Body_x[2986];
                c_Body_y[2986] = n_Body_y[2986];
                c_Body_x[2987] = n_Body_x[2987];
                c_Body_y[2987] = n_Body_y[2987];
                c_Body_x[2988] = n_Body_x[2988];
                c_Body_y[2988] = n_Body_y[2988];
                c_Body_x[2989] = n_Body_x[2989];
                c_Body_y[2989] = n_Body_y[2989];
                c_Body_x[2990] = n_Body_x[2990];
                c_Body_y[2990] = n_Body_y[2990];
                c_Body_x[2991] = n_Body_x[2991];
                c_Body_y[2991] = n_Body_y[2991];
                c_Body_x[2992] = n_Body_x[2992];
                c_Body_y[2992] = n_Body_y[2992];
                c_Body_x[2993] = n_Body_x[2993];
                c_Body_y[2993] = n_Body_y[2993];
                c_Body_x[2994] = n_Body_x[2994];
                c_Body_y[2994] = n_Body_y[2994];
                c_Body_x[2995] = n_Body_x[2995];
                c_Body_y[2995] = n_Body_y[2995];
                c_Body_x[2996] = n_Body_x[2996];
                c_Body_y[2996] = n_Body_y[2996];
                c_Body_x[2997] = n_Body_x[2997];
                c_Body_y[2997] = n_Body_y[2997];
                c_Body_x[2998] = n_Body_x[2998];
                c_Body_y[2998] = n_Body_y[2998];
                c_Body_x[2999] = n_Body_x[2999];
                c_Body_y[2999] = n_Body_y[2999];
                c_Body_x[3000] = n_Body_x[3000];
                c_Body_y[3000] = n_Body_y[3000];
                c_Body_x[3001] = n_Body_x[3001];
                c_Body_y[3001] = n_Body_y[3001];
                c_Body_x[3002] = n_Body_x[3002];
                c_Body_y[3002] = n_Body_y[3002];
                c_Body_x[3003] = n_Body_x[3003];
                c_Body_y[3003] = n_Body_y[3003];
                c_Body_x[3004] = n_Body_x[3004];
                c_Body_y[3004] = n_Body_y[3004];
                c_Body_x[3005] = n_Body_x[3005];
                c_Body_y[3005] = n_Body_y[3005];
                c_Body_x[3006] = n_Body_x[3006];
                c_Body_y[3006] = n_Body_y[3006];
                c_Body_x[3007] = n_Body_x[3007];
                c_Body_y[3007] = n_Body_y[3007];
                c_Body_x[3008] = n_Body_x[3008];
                c_Body_y[3008] = n_Body_y[3008];
                c_Body_x[3009] = n_Body_x[3009];
                c_Body_y[3009] = n_Body_y[3009];
                c_Body_x[3010] = n_Body_x[3010];
                c_Body_y[3010] = n_Body_y[3010];
                c_Body_x[3011] = n_Body_x[3011];
                c_Body_y[3011] = n_Body_y[3011];
                c_Body_x[3012] = n_Body_x[3012];
                c_Body_y[3012] = n_Body_y[3012];
                c_Body_x[3013] = n_Body_x[3013];
                c_Body_y[3013] = n_Body_y[3013];
                c_Body_x[3014] = n_Body_x[3014];
                c_Body_y[3014] = n_Body_y[3014];
                c_Body_x[3015] = n_Body_x[3015];
                c_Body_y[3015] = n_Body_y[3015];
                c_Body_x[3016] = n_Body_x[3016];
                c_Body_y[3016] = n_Body_y[3016];
                c_Body_x[3017] = n_Body_x[3017];
                c_Body_y[3017] = n_Body_y[3017];
                c_Body_x[3018] = n_Body_x[3018];
                c_Body_y[3018] = n_Body_y[3018];
                c_Body_x[3019] = n_Body_x[3019];
                c_Body_y[3019] = n_Body_y[3019];
                c_Body_x[3020] = n_Body_x[3020];
                c_Body_y[3020] = n_Body_y[3020];
                c_Body_x[3021] = n_Body_x[3021];
                c_Body_y[3021] = n_Body_y[3021];
                c_Body_x[3022] = n_Body_x[3022];
                c_Body_y[3022] = n_Body_y[3022];
                c_Body_x[3023] = n_Body_x[3023];
                c_Body_y[3023] = n_Body_y[3023];
                c_Body_x[3024] = n_Body_x[3024];
                c_Body_y[3024] = n_Body_y[3024];
                c_Body_x[3025] = n_Body_x[3025];
                c_Body_y[3025] = n_Body_y[3025];
                c_Body_x[3026] = n_Body_x[3026];
                c_Body_y[3026] = n_Body_y[3026];
                c_Body_x[3027] = n_Body_x[3027];
                c_Body_y[3027] = n_Body_y[3027];
                c_Body_x[3028] = n_Body_x[3028];
                c_Body_y[3028] = n_Body_y[3028];
                c_Body_x[3029] = n_Body_x[3029];
                c_Body_y[3029] = n_Body_y[3029];
                c_Body_x[3030] = n_Body_x[3030];
                c_Body_y[3030] = n_Body_y[3030];
                c_Body_x[3031] = n_Body_x[3031];
                c_Body_y[3031] = n_Body_y[3031];
                c_Body_x[3032] = n_Body_x[3032];
                c_Body_y[3032] = n_Body_y[3032];
                c_Body_x[3033] = n_Body_x[3033];
                c_Body_y[3033] = n_Body_y[3033];
                c_Body_x[3034] = n_Body_x[3034];
                c_Body_y[3034] = n_Body_y[3034];
                c_Body_x[3035] = n_Body_x[3035];
                c_Body_y[3035] = n_Body_y[3035];
                c_Body_x[3036] = n_Body_x[3036];
                c_Body_y[3036] = n_Body_y[3036];
                c_Body_x[3037] = n_Body_x[3037];
                c_Body_y[3037] = n_Body_y[3037];
                c_Body_x[3038] = n_Body_x[3038];
                c_Body_y[3038] = n_Body_y[3038];
                c_Body_x[3039] = n_Body_x[3039];
                c_Body_y[3039] = n_Body_y[3039];
                c_Body_x[3040] = n_Body_x[3040];
                c_Body_y[3040] = n_Body_y[3040];
                c_Body_x[3041] = n_Body_x[3041];
                c_Body_y[3041] = n_Body_y[3041];
                c_Body_x[3042] = n_Body_x[3042];
                c_Body_y[3042] = n_Body_y[3042];
                c_Body_x[3043] = n_Body_x[3043];
                c_Body_y[3043] = n_Body_y[3043];
                c_Body_x[3044] = n_Body_x[3044];
                c_Body_y[3044] = n_Body_y[3044];
                c_Body_x[3045] = n_Body_x[3045];
                c_Body_y[3045] = n_Body_y[3045];
                c_Body_x[3046] = n_Body_x[3046];
                c_Body_y[3046] = n_Body_y[3046];
                c_Body_x[3047] = n_Body_x[3047];
                c_Body_y[3047] = n_Body_y[3047];
                c_Body_x[3048] = n_Body_x[3048];
                c_Body_y[3048] = n_Body_y[3048];
                c_Body_x[3049] = n_Body_x[3049];
                c_Body_y[3049] = n_Body_y[3049];
                c_Body_x[3050] = n_Body_x[3050];
                c_Body_y[3050] = n_Body_y[3050];
                c_Body_x[3051] = n_Body_x[3051];
                c_Body_y[3051] = n_Body_y[3051];
                c_Body_x[3052] = n_Body_x[3052];
                c_Body_y[3052] = n_Body_y[3052];
                c_Body_x[3053] = n_Body_x[3053];
                c_Body_y[3053] = n_Body_y[3053];
                c_Body_x[3054] = n_Body_x[3054];
                c_Body_y[3054] = n_Body_y[3054];
                c_Body_x[3055] = n_Body_x[3055];
                c_Body_y[3055] = n_Body_y[3055];
                c_Body_x[3056] = n_Body_x[3056];
                c_Body_y[3056] = n_Body_y[3056];
                c_Body_x[3057] = n_Body_x[3057];
                c_Body_y[3057] = n_Body_y[3057];
                c_Body_x[3058] = n_Body_x[3058];
                c_Body_y[3058] = n_Body_y[3058];
                c_Body_x[3059] = n_Body_x[3059];
                c_Body_y[3059] = n_Body_y[3059];
                c_Body_x[3060] = n_Body_x[3060];
                c_Body_y[3060] = n_Body_y[3060];
                c_Body_x[3061] = n_Body_x[3061];
                c_Body_y[3061] = n_Body_y[3061];
                c_Body_x[3062] = n_Body_x[3062];
                c_Body_y[3062] = n_Body_y[3062];
                c_Body_x[3063] = n_Body_x[3063];
                c_Body_y[3063] = n_Body_y[3063];
                c_Body_x[3064] = n_Body_x[3064];
                c_Body_y[3064] = n_Body_y[3064];
                c_Body_x[3065] = n_Body_x[3065];
                c_Body_y[3065] = n_Body_y[3065];
                c_Body_x[3066] = n_Body_x[3066];
                c_Body_y[3066] = n_Body_y[3066];
                c_Body_x[3067] = n_Body_x[3067];
                c_Body_y[3067] = n_Body_y[3067];
                c_Body_x[3068] = n_Body_x[3068];
                c_Body_y[3068] = n_Body_y[3068];
                c_Body_x[3069] = n_Body_x[3069];
                c_Body_y[3069] = n_Body_y[3069];
                c_Body_x[3070] = n_Body_x[3070];
                c_Body_y[3070] = n_Body_y[3070];
                c_Body_x[3071] = n_Body_x[3071];
                c_Body_y[3071] = n_Body_y[3071];

        end
    end

    // SetHead모듈 연결
    SetHead SH0 (i_Clk, i_Rst,
                 c_Way, c_Push, c_Head_x, c_Head_y,
                 SH_o_Head_x, SH_o_Head_y, SH_o_Way);

    // 점수, 속도 모듈 연결
    wire [3:0] SF_o_F0, SF_o_F1, CF_o_F0, CF_o_F1, CF_o_F2, CF_o_F3;
    SpeedFND SF0(c_Speed, SF_o_F0, SF_o_F1);
    ScoreFND CF0(c_Size, CF_o_F0, CF_o_F1, CF_o_F2, CF_o_F3);
    FND F0(SF_o_F0, o_Speed_FND0);
    FND F1(SF_o_F1, o_Speed_FND1);
    FND F2(CF_o_F0, o_Score_FND0);
    FND F3(CF_o_F0, o_Score_FND1);
    FND F4(CF_o_F0, o_Score_FND2);
    FND F5(CF_o_F0, o_Score_FND3);

    //VGA모듈 연결
    output o_hsync, o_vsync;
    output [7:0] o_red, o_green, o_blue;
    Vga V0(i_Clk, i_Rst, i_Body_x_flat, i_Body_y_flat, c_Item_x, c_Item_y, c_Size,
           o_hsync, o_vsync, o_red, o_blue, o_green);

    wire o_isMakeItem_Done;

    always @* begin
        n_Head_x = c_Head_x;
        n_Head_y = c_Head_y;
        n_Item_x = c_Item_x;
        n_Item_y = c_Item_y;
        n_Size   = c_Size;
        n_ClkCnt = 0;
        n_Way    = c_Way;
        n_Push   = c_Push;
        n_State  = c_State;
        n_Speed  = c_Speed;
        n_SpdTimeCnt = c_SpdTimeCnt;
        
        //무수히 많은 대입문들...
            n_Body_x[0] = c_Body_x[0];
            n_Body_y[0] = c_Body_y[0];
            n_Body_x[1] = c_Body_x[1];
            n_Body_y[1] = c_Body_y[1];
            n_Body_x[2] = c_Body_x[2];
            n_Body_y[2] = c_Body_y[2];
            n_Body_x[3] = c_Body_x[3];
            n_Body_y[3] = c_Body_y[3];
            n_Body_x[4] = c_Body_x[4];
            n_Body_y[4] = c_Body_y[4];
            n_Body_x[5] = c_Body_x[5];
            n_Body_y[5] = c_Body_y[5];
            n_Body_x[6] = c_Body_x[6];
            n_Body_y[6] = c_Body_y[6];
            n_Body_x[7] = c_Body_x[7];
            n_Body_y[7] = c_Body_y[7];
            n_Body_x[8] = c_Body_x[8];
            n_Body_y[8] = c_Body_y[8];
            n_Body_x[9] = c_Body_x[9];
            n_Body_y[9] = c_Body_y[9];
            n_Body_x[10] = c_Body_x[10];
            n_Body_y[10] = c_Body_y[10];
            n_Body_x[11] = c_Body_x[11];
            n_Body_y[11] = c_Body_y[11];
            n_Body_x[12] = c_Body_x[12];
            n_Body_y[12] = c_Body_y[12];
            n_Body_x[13] = c_Body_x[13];
            n_Body_y[13] = c_Body_y[13];
            n_Body_x[14] = c_Body_x[14];
            n_Body_y[14] = c_Body_y[14];
            n_Body_x[15] = c_Body_x[15];
            n_Body_y[15] = c_Body_y[15];
            n_Body_x[16] = c_Body_x[16];
            n_Body_y[16] = c_Body_y[16];
            n_Body_x[17] = c_Body_x[17];
            n_Body_y[17] = c_Body_y[17];
            n_Body_x[18] = c_Body_x[18];
            n_Body_y[18] = c_Body_y[18];
            n_Body_x[19] = c_Body_x[19];
            n_Body_y[19] = c_Body_y[19];
            n_Body_x[20] = c_Body_x[20];
            n_Body_y[20] = c_Body_y[20];
            n_Body_x[21] = c_Body_x[21];
            n_Body_y[21] = c_Body_y[21];
            n_Body_x[22] = c_Body_x[22];
            n_Body_y[22] = c_Body_y[22];
            n_Body_x[23] = c_Body_x[23];
            n_Body_y[23] = c_Body_y[23];
            n_Body_x[24] = c_Body_x[24];
            n_Body_y[24] = c_Body_y[24];
            n_Body_x[25] = c_Body_x[25];
            n_Body_y[25] = c_Body_y[25];
            n_Body_x[26] = c_Body_x[26];
            n_Body_y[26] = c_Body_y[26];
            n_Body_x[27] = c_Body_x[27];
            n_Body_y[27] = c_Body_y[27];
            n_Body_x[28] = c_Body_x[28];
            n_Body_y[28] = c_Body_y[28];
            n_Body_x[29] = c_Body_x[29];
            n_Body_y[29] = c_Body_y[29];
            n_Body_x[30] = c_Body_x[30];
            n_Body_y[30] = c_Body_y[30];
            n_Body_x[31] = c_Body_x[31];
            n_Body_y[31] = c_Body_y[31];
            n_Body_x[32] = c_Body_x[32];
            n_Body_y[32] = c_Body_y[32];
            n_Body_x[33] = c_Body_x[33];
            n_Body_y[33] = c_Body_y[33];
            n_Body_x[34] = c_Body_x[34];
            n_Body_y[34] = c_Body_y[34];
            n_Body_x[35] = c_Body_x[35];
            n_Body_y[35] = c_Body_y[35];
            n_Body_x[36] = c_Body_x[36];
            n_Body_y[36] = c_Body_y[36];
            n_Body_x[37] = c_Body_x[37];
            n_Body_y[37] = c_Body_y[37];
            n_Body_x[38] = c_Body_x[38];
            n_Body_y[38] = c_Body_y[38];
            n_Body_x[39] = c_Body_x[39];
            n_Body_y[39] = c_Body_y[39];
            n_Body_x[40] = c_Body_x[40];
            n_Body_y[40] = c_Body_y[40];
            n_Body_x[41] = c_Body_x[41];
            n_Body_y[41] = c_Body_y[41];
            n_Body_x[42] = c_Body_x[42];
            n_Body_y[42] = c_Body_y[42];
            n_Body_x[43] = c_Body_x[43];
            n_Body_y[43] = c_Body_y[43];
            n_Body_x[44] = c_Body_x[44];
            n_Body_y[44] = c_Body_y[44];
            n_Body_x[45] = c_Body_x[45];
            n_Body_y[45] = c_Body_y[45];
            n_Body_x[46] = c_Body_x[46];
            n_Body_y[46] = c_Body_y[46];
            n_Body_x[47] = c_Body_x[47];
            n_Body_y[47] = c_Body_y[47];
            n_Body_x[48] = c_Body_x[48];
            n_Body_y[48] = c_Body_y[48];
            n_Body_x[49] = c_Body_x[49];
            n_Body_y[49] = c_Body_y[49];
            n_Body_x[50] = c_Body_x[50];
            n_Body_y[50] = c_Body_y[50];
            n_Body_x[51] = c_Body_x[51];
            n_Body_y[51] = c_Body_y[51];
            n_Body_x[52] = c_Body_x[52];
            n_Body_y[52] = c_Body_y[52];
            n_Body_x[53] = c_Body_x[53];
            n_Body_y[53] = c_Body_y[53];
            n_Body_x[54] = c_Body_x[54];
            n_Body_y[54] = c_Body_y[54];
            n_Body_x[55] = c_Body_x[55];
            n_Body_y[55] = c_Body_y[55];
            n_Body_x[56] = c_Body_x[56];
            n_Body_y[56] = c_Body_y[56];
            n_Body_x[57] = c_Body_x[57];
            n_Body_y[57] = c_Body_y[57];
            n_Body_x[58] = c_Body_x[58];
            n_Body_y[58] = c_Body_y[58];
            n_Body_x[59] = c_Body_x[59];
            n_Body_y[59] = c_Body_y[59];
            n_Body_x[60] = c_Body_x[60];
            n_Body_y[60] = c_Body_y[60];
            n_Body_x[61] = c_Body_x[61];
            n_Body_y[61] = c_Body_y[61];
            n_Body_x[62] = c_Body_x[62];
            n_Body_y[62] = c_Body_y[62];
            n_Body_x[63] = c_Body_x[63];
            n_Body_y[63] = c_Body_y[63];
            n_Body_x[64] = c_Body_x[64];
            n_Body_y[64] = c_Body_y[64];
            n_Body_x[65] = c_Body_x[65];
            n_Body_y[65] = c_Body_y[65];
            n_Body_x[66] = c_Body_x[66];
            n_Body_y[66] = c_Body_y[66];
            n_Body_x[67] = c_Body_x[67];
            n_Body_y[67] = c_Body_y[67];
            n_Body_x[68] = c_Body_x[68];
            n_Body_y[68] = c_Body_y[68];
            n_Body_x[69] = c_Body_x[69];
            n_Body_y[69] = c_Body_y[69];
            n_Body_x[70] = c_Body_x[70];
            n_Body_y[70] = c_Body_y[70];
            n_Body_x[71] = c_Body_x[71];
            n_Body_y[71] = c_Body_y[71];
            n_Body_x[72] = c_Body_x[72];
            n_Body_y[72] = c_Body_y[72];
            n_Body_x[73] = c_Body_x[73];
            n_Body_y[73] = c_Body_y[73];
            n_Body_x[74] = c_Body_x[74];
            n_Body_y[74] = c_Body_y[74];
            n_Body_x[75] = c_Body_x[75];
            n_Body_y[75] = c_Body_y[75];
            n_Body_x[76] = c_Body_x[76];
            n_Body_y[76] = c_Body_y[76];
            n_Body_x[77] = c_Body_x[77];
            n_Body_y[77] = c_Body_y[77];
            n_Body_x[78] = c_Body_x[78];
            n_Body_y[78] = c_Body_y[78];
            n_Body_x[79] = c_Body_x[79];
            n_Body_y[79] = c_Body_y[79];
            n_Body_x[80] = c_Body_x[80];
            n_Body_y[80] = c_Body_y[80];
            n_Body_x[81] = c_Body_x[81];
            n_Body_y[81] = c_Body_y[81];
            n_Body_x[82] = c_Body_x[82];
            n_Body_y[82] = c_Body_y[82];
            n_Body_x[83] = c_Body_x[83];
            n_Body_y[83] = c_Body_y[83];
            n_Body_x[84] = c_Body_x[84];
            n_Body_y[84] = c_Body_y[84];
            n_Body_x[85] = c_Body_x[85];
            n_Body_y[85] = c_Body_y[85];
            n_Body_x[86] = c_Body_x[86];
            n_Body_y[86] = c_Body_y[86];
            n_Body_x[87] = c_Body_x[87];
            n_Body_y[87] = c_Body_y[87];
            n_Body_x[88] = c_Body_x[88];
            n_Body_y[88] = c_Body_y[88];
            n_Body_x[89] = c_Body_x[89];
            n_Body_y[89] = c_Body_y[89];
            n_Body_x[90] = c_Body_x[90];
            n_Body_y[90] = c_Body_y[90];
            n_Body_x[91] = c_Body_x[91];
            n_Body_y[91] = c_Body_y[91];
            n_Body_x[92] = c_Body_x[92];
            n_Body_y[92] = c_Body_y[92];
            n_Body_x[93] = c_Body_x[93];
            n_Body_y[93] = c_Body_y[93];
            n_Body_x[94] = c_Body_x[94];
            n_Body_y[94] = c_Body_y[94];
            n_Body_x[95] = c_Body_x[95];
            n_Body_y[95] = c_Body_y[95];
            n_Body_x[96] = c_Body_x[96];
            n_Body_y[96] = c_Body_y[96];
            n_Body_x[97] = c_Body_x[97];
            n_Body_y[97] = c_Body_y[97];
            n_Body_x[98] = c_Body_x[98];
            n_Body_y[98] = c_Body_y[98];
            n_Body_x[99] = c_Body_x[99];
            n_Body_y[99] = c_Body_y[99];
            n_Body_x[100] = c_Body_x[100];
            n_Body_y[100] = c_Body_y[100];
            n_Body_x[101] = c_Body_x[101];
            n_Body_y[101] = c_Body_y[101];
            n_Body_x[102] = c_Body_x[102];
            n_Body_y[102] = c_Body_y[102];
            n_Body_x[103] = c_Body_x[103];
            n_Body_y[103] = c_Body_y[103];
            n_Body_x[104] = c_Body_x[104];
            n_Body_y[104] = c_Body_y[104];
            n_Body_x[105] = c_Body_x[105];
            n_Body_y[105] = c_Body_y[105];
            n_Body_x[106] = c_Body_x[106];
            n_Body_y[106] = c_Body_y[106];
            n_Body_x[107] = c_Body_x[107];
            n_Body_y[107] = c_Body_y[107];
            n_Body_x[108] = c_Body_x[108];
            n_Body_y[108] = c_Body_y[108];
            n_Body_x[109] = c_Body_x[109];
            n_Body_y[109] = c_Body_y[109];
            n_Body_x[110] = c_Body_x[110];
            n_Body_y[110] = c_Body_y[110];
            n_Body_x[111] = c_Body_x[111];
            n_Body_y[111] = c_Body_y[111];
            n_Body_x[112] = c_Body_x[112];
            n_Body_y[112] = c_Body_y[112];
            n_Body_x[113] = c_Body_x[113];
            n_Body_y[113] = c_Body_y[113];
            n_Body_x[114] = c_Body_x[114];
            n_Body_y[114] = c_Body_y[114];
            n_Body_x[115] = c_Body_x[115];
            n_Body_y[115] = c_Body_y[115];
            n_Body_x[116] = c_Body_x[116];
            n_Body_y[116] = c_Body_y[116];
            n_Body_x[117] = c_Body_x[117];
            n_Body_y[117] = c_Body_y[117];
            n_Body_x[118] = c_Body_x[118];
            n_Body_y[118] = c_Body_y[118];
            n_Body_x[119] = c_Body_x[119];
            n_Body_y[119] = c_Body_y[119];
            n_Body_x[120] = c_Body_x[120];
            n_Body_y[120] = c_Body_y[120];
            n_Body_x[121] = c_Body_x[121];
            n_Body_y[121] = c_Body_y[121];
            n_Body_x[122] = c_Body_x[122];
            n_Body_y[122] = c_Body_y[122];
            n_Body_x[123] = c_Body_x[123];
            n_Body_y[123] = c_Body_y[123];
            n_Body_x[124] = c_Body_x[124];
            n_Body_y[124] = c_Body_y[124];
            n_Body_x[125] = c_Body_x[125];
            n_Body_y[125] = c_Body_y[125];
            n_Body_x[126] = c_Body_x[126];
            n_Body_y[126] = c_Body_y[126];
            n_Body_x[127] = c_Body_x[127];
            n_Body_y[127] = c_Body_y[127];
            n_Body_x[128] = c_Body_x[128];
            n_Body_y[128] = c_Body_y[128];
            n_Body_x[129] = c_Body_x[129];
            n_Body_y[129] = c_Body_y[129];
            n_Body_x[130] = c_Body_x[130];
            n_Body_y[130] = c_Body_y[130];
            n_Body_x[131] = c_Body_x[131];
            n_Body_y[131] = c_Body_y[131];
            n_Body_x[132] = c_Body_x[132];
            n_Body_y[132] = c_Body_y[132];
            n_Body_x[133] = c_Body_x[133];
            n_Body_y[133] = c_Body_y[133];
            n_Body_x[134] = c_Body_x[134];
            n_Body_y[134] = c_Body_y[134];
            n_Body_x[135] = c_Body_x[135];
            n_Body_y[135] = c_Body_y[135];
            n_Body_x[136] = c_Body_x[136];
            n_Body_y[136] = c_Body_y[136];
            n_Body_x[137] = c_Body_x[137];
            n_Body_y[137] = c_Body_y[137];
            n_Body_x[138] = c_Body_x[138];
            n_Body_y[138] = c_Body_y[138];
            n_Body_x[139] = c_Body_x[139];
            n_Body_y[139] = c_Body_y[139];
            n_Body_x[140] = c_Body_x[140];
            n_Body_y[140] = c_Body_y[140];
            n_Body_x[141] = c_Body_x[141];
            n_Body_y[141] = c_Body_y[141];
            n_Body_x[142] = c_Body_x[142];
            n_Body_y[142] = c_Body_y[142];
            n_Body_x[143] = c_Body_x[143];
            n_Body_y[143] = c_Body_y[143];
            n_Body_x[144] = c_Body_x[144];
            n_Body_y[144] = c_Body_y[144];
            n_Body_x[145] = c_Body_x[145];
            n_Body_y[145] = c_Body_y[145];
            n_Body_x[146] = c_Body_x[146];
            n_Body_y[146] = c_Body_y[146];
            n_Body_x[147] = c_Body_x[147];
            n_Body_y[147] = c_Body_y[147];
            n_Body_x[148] = c_Body_x[148];
            n_Body_y[148] = c_Body_y[148];
            n_Body_x[149] = c_Body_x[149];
            n_Body_y[149] = c_Body_y[149];
            n_Body_x[150] = c_Body_x[150];
            n_Body_y[150] = c_Body_y[150];
            n_Body_x[151] = c_Body_x[151];
            n_Body_y[151] = c_Body_y[151];
            n_Body_x[152] = c_Body_x[152];
            n_Body_y[152] = c_Body_y[152];
            n_Body_x[153] = c_Body_x[153];
            n_Body_y[153] = c_Body_y[153];
            n_Body_x[154] = c_Body_x[154];
            n_Body_y[154] = c_Body_y[154];
            n_Body_x[155] = c_Body_x[155];
            n_Body_y[155] = c_Body_y[155];
            n_Body_x[156] = c_Body_x[156];
            n_Body_y[156] = c_Body_y[156];
            n_Body_x[157] = c_Body_x[157];
            n_Body_y[157] = c_Body_y[157];
            n_Body_x[158] = c_Body_x[158];
            n_Body_y[158] = c_Body_y[158];
            n_Body_x[159] = c_Body_x[159];
            n_Body_y[159] = c_Body_y[159];
            n_Body_x[160] = c_Body_x[160];
            n_Body_y[160] = c_Body_y[160];
            n_Body_x[161] = c_Body_x[161];
            n_Body_y[161] = c_Body_y[161];
            n_Body_x[162] = c_Body_x[162];
            n_Body_y[162] = c_Body_y[162];
            n_Body_x[163] = c_Body_x[163];
            n_Body_y[163] = c_Body_y[163];
            n_Body_x[164] = c_Body_x[164];
            n_Body_y[164] = c_Body_y[164];
            n_Body_x[165] = c_Body_x[165];
            n_Body_y[165] = c_Body_y[165];
            n_Body_x[166] = c_Body_x[166];
            n_Body_y[166] = c_Body_y[166];
            n_Body_x[167] = c_Body_x[167];
            n_Body_y[167] = c_Body_y[167];
            n_Body_x[168] = c_Body_x[168];
            n_Body_y[168] = c_Body_y[168];
            n_Body_x[169] = c_Body_x[169];
            n_Body_y[169] = c_Body_y[169];
            n_Body_x[170] = c_Body_x[170];
            n_Body_y[170] = c_Body_y[170];
            n_Body_x[171] = c_Body_x[171];
            n_Body_y[171] = c_Body_y[171];
            n_Body_x[172] = c_Body_x[172];
            n_Body_y[172] = c_Body_y[172];
            n_Body_x[173] = c_Body_x[173];
            n_Body_y[173] = c_Body_y[173];
            n_Body_x[174] = c_Body_x[174];
            n_Body_y[174] = c_Body_y[174];
            n_Body_x[175] = c_Body_x[175];
            n_Body_y[175] = c_Body_y[175];
            n_Body_x[176] = c_Body_x[176];
            n_Body_y[176] = c_Body_y[176];
            n_Body_x[177] = c_Body_x[177];
            n_Body_y[177] = c_Body_y[177];
            n_Body_x[178] = c_Body_x[178];
            n_Body_y[178] = c_Body_y[178];
            n_Body_x[179] = c_Body_x[179];
            n_Body_y[179] = c_Body_y[179];
            n_Body_x[180] = c_Body_x[180];
            n_Body_y[180] = c_Body_y[180];
            n_Body_x[181] = c_Body_x[181];
            n_Body_y[181] = c_Body_y[181];
            n_Body_x[182] = c_Body_x[182];
            n_Body_y[182] = c_Body_y[182];
            n_Body_x[183] = c_Body_x[183];
            n_Body_y[183] = c_Body_y[183];
            n_Body_x[184] = c_Body_x[184];
            n_Body_y[184] = c_Body_y[184];
            n_Body_x[185] = c_Body_x[185];
            n_Body_y[185] = c_Body_y[185];
            n_Body_x[186] = c_Body_x[186];
            n_Body_y[186] = c_Body_y[186];
            n_Body_x[187] = c_Body_x[187];
            n_Body_y[187] = c_Body_y[187];
            n_Body_x[188] = c_Body_x[188];
            n_Body_y[188] = c_Body_y[188];
            n_Body_x[189] = c_Body_x[189];
            n_Body_y[189] = c_Body_y[189];
            n_Body_x[190] = c_Body_x[190];
            n_Body_y[190] = c_Body_y[190];
            n_Body_x[191] = c_Body_x[191];
            n_Body_y[191] = c_Body_y[191];
            n_Body_x[192] = c_Body_x[192];
            n_Body_y[192] = c_Body_y[192];
            n_Body_x[193] = c_Body_x[193];
            n_Body_y[193] = c_Body_y[193];
            n_Body_x[194] = c_Body_x[194];
            n_Body_y[194] = c_Body_y[194];
            n_Body_x[195] = c_Body_x[195];
            n_Body_y[195] = c_Body_y[195];
            n_Body_x[196] = c_Body_x[196];
            n_Body_y[196] = c_Body_y[196];
            n_Body_x[197] = c_Body_x[197];
            n_Body_y[197] = c_Body_y[197];
            n_Body_x[198] = c_Body_x[198];
            n_Body_y[198] = c_Body_y[198];
            n_Body_x[199] = c_Body_x[199];
            n_Body_y[199] = c_Body_y[199];
            n_Body_x[200] = c_Body_x[200];
            n_Body_y[200] = c_Body_y[200];
            n_Body_x[201] = c_Body_x[201];
            n_Body_y[201] = c_Body_y[201];
            n_Body_x[202] = c_Body_x[202];
            n_Body_y[202] = c_Body_y[202];
            n_Body_x[203] = c_Body_x[203];
            n_Body_y[203] = c_Body_y[203];
            n_Body_x[204] = c_Body_x[204];
            n_Body_y[204] = c_Body_y[204];
            n_Body_x[205] = c_Body_x[205];
            n_Body_y[205] = c_Body_y[205];
            n_Body_x[206] = c_Body_x[206];
            n_Body_y[206] = c_Body_y[206];
            n_Body_x[207] = c_Body_x[207];
            n_Body_y[207] = c_Body_y[207];
            n_Body_x[208] = c_Body_x[208];
            n_Body_y[208] = c_Body_y[208];
            n_Body_x[209] = c_Body_x[209];
            n_Body_y[209] = c_Body_y[209];
            n_Body_x[210] = c_Body_x[210];
            n_Body_y[210] = c_Body_y[210];
            n_Body_x[211] = c_Body_x[211];
            n_Body_y[211] = c_Body_y[211];
            n_Body_x[212] = c_Body_x[212];
            n_Body_y[212] = c_Body_y[212];
            n_Body_x[213] = c_Body_x[213];
            n_Body_y[213] = c_Body_y[213];
            n_Body_x[214] = c_Body_x[214];
            n_Body_y[214] = c_Body_y[214];
            n_Body_x[215] = c_Body_x[215];
            n_Body_y[215] = c_Body_y[215];
            n_Body_x[216] = c_Body_x[216];
            n_Body_y[216] = c_Body_y[216];
            n_Body_x[217] = c_Body_x[217];
            n_Body_y[217] = c_Body_y[217];
            n_Body_x[218] = c_Body_x[218];
            n_Body_y[218] = c_Body_y[218];
            n_Body_x[219] = c_Body_x[219];
            n_Body_y[219] = c_Body_y[219];
            n_Body_x[220] = c_Body_x[220];
            n_Body_y[220] = c_Body_y[220];
            n_Body_x[221] = c_Body_x[221];
            n_Body_y[221] = c_Body_y[221];
            n_Body_x[222] = c_Body_x[222];
            n_Body_y[222] = c_Body_y[222];
            n_Body_x[223] = c_Body_x[223];
            n_Body_y[223] = c_Body_y[223];
            n_Body_x[224] = c_Body_x[224];
            n_Body_y[224] = c_Body_y[224];
            n_Body_x[225] = c_Body_x[225];
            n_Body_y[225] = c_Body_y[225];
            n_Body_x[226] = c_Body_x[226];
            n_Body_y[226] = c_Body_y[226];
            n_Body_x[227] = c_Body_x[227];
            n_Body_y[227] = c_Body_y[227];
            n_Body_x[228] = c_Body_x[228];
            n_Body_y[228] = c_Body_y[228];
            n_Body_x[229] = c_Body_x[229];
            n_Body_y[229] = c_Body_y[229];
            n_Body_x[230] = c_Body_x[230];
            n_Body_y[230] = c_Body_y[230];
            n_Body_x[231] = c_Body_x[231];
            n_Body_y[231] = c_Body_y[231];
            n_Body_x[232] = c_Body_x[232];
            n_Body_y[232] = c_Body_y[232];
            n_Body_x[233] = c_Body_x[233];
            n_Body_y[233] = c_Body_y[233];
            n_Body_x[234] = c_Body_x[234];
            n_Body_y[234] = c_Body_y[234];
            n_Body_x[235] = c_Body_x[235];
            n_Body_y[235] = c_Body_y[235];
            n_Body_x[236] = c_Body_x[236];
            n_Body_y[236] = c_Body_y[236];
            n_Body_x[237] = c_Body_x[237];
            n_Body_y[237] = c_Body_y[237];
            n_Body_x[238] = c_Body_x[238];
            n_Body_y[238] = c_Body_y[238];
            n_Body_x[239] = c_Body_x[239];
            n_Body_y[239] = c_Body_y[239];
            n_Body_x[240] = c_Body_x[240];
            n_Body_y[240] = c_Body_y[240];
            n_Body_x[241] = c_Body_x[241];
            n_Body_y[241] = c_Body_y[241];
            n_Body_x[242] = c_Body_x[242];
            n_Body_y[242] = c_Body_y[242];
            n_Body_x[243] = c_Body_x[243];
            n_Body_y[243] = c_Body_y[243];
            n_Body_x[244] = c_Body_x[244];
            n_Body_y[244] = c_Body_y[244];
            n_Body_x[245] = c_Body_x[245];
            n_Body_y[245] = c_Body_y[245];
            n_Body_x[246] = c_Body_x[246];
            n_Body_y[246] = c_Body_y[246];
            n_Body_x[247] = c_Body_x[247];
            n_Body_y[247] = c_Body_y[247];
            n_Body_x[248] = c_Body_x[248];
            n_Body_y[248] = c_Body_y[248];
            n_Body_x[249] = c_Body_x[249];
            n_Body_y[249] = c_Body_y[249];
            n_Body_x[250] = c_Body_x[250];
            n_Body_y[250] = c_Body_y[250];
            n_Body_x[251] = c_Body_x[251];
            n_Body_y[251] = c_Body_y[251];
            n_Body_x[252] = c_Body_x[252];
            n_Body_y[252] = c_Body_y[252];
            n_Body_x[253] = c_Body_x[253];
            n_Body_y[253] = c_Body_y[253];
            n_Body_x[254] = c_Body_x[254];
            n_Body_y[254] = c_Body_y[254];
            n_Body_x[255] = c_Body_x[255];
            n_Body_y[255] = c_Body_y[255];
            n_Body_x[256] = c_Body_x[256];
            n_Body_y[256] = c_Body_y[256];
            n_Body_x[257] = c_Body_x[257];
            n_Body_y[257] = c_Body_y[257];
            n_Body_x[258] = c_Body_x[258];
            n_Body_y[258] = c_Body_y[258];
            n_Body_x[259] = c_Body_x[259];
            n_Body_y[259] = c_Body_y[259];
            n_Body_x[260] = c_Body_x[260];
            n_Body_y[260] = c_Body_y[260];
            n_Body_x[261] = c_Body_x[261];
            n_Body_y[261] = c_Body_y[261];
            n_Body_x[262] = c_Body_x[262];
            n_Body_y[262] = c_Body_y[262];
            n_Body_x[263] = c_Body_x[263];
            n_Body_y[263] = c_Body_y[263];
            n_Body_x[264] = c_Body_x[264];
            n_Body_y[264] = c_Body_y[264];
            n_Body_x[265] = c_Body_x[265];
            n_Body_y[265] = c_Body_y[265];
            n_Body_x[266] = c_Body_x[266];
            n_Body_y[266] = c_Body_y[266];
            n_Body_x[267] = c_Body_x[267];
            n_Body_y[267] = c_Body_y[267];
            n_Body_x[268] = c_Body_x[268];
            n_Body_y[268] = c_Body_y[268];
            n_Body_x[269] = c_Body_x[269];
            n_Body_y[269] = c_Body_y[269];
            n_Body_x[270] = c_Body_x[270];
            n_Body_y[270] = c_Body_y[270];
            n_Body_x[271] = c_Body_x[271];
            n_Body_y[271] = c_Body_y[271];
            n_Body_x[272] = c_Body_x[272];
            n_Body_y[272] = c_Body_y[272];
            n_Body_x[273] = c_Body_x[273];
            n_Body_y[273] = c_Body_y[273];
            n_Body_x[274] = c_Body_x[274];
            n_Body_y[274] = c_Body_y[274];
            n_Body_x[275] = c_Body_x[275];
            n_Body_y[275] = c_Body_y[275];
            n_Body_x[276] = c_Body_x[276];
            n_Body_y[276] = c_Body_y[276];
            n_Body_x[277] = c_Body_x[277];
            n_Body_y[277] = c_Body_y[277];
            n_Body_x[278] = c_Body_x[278];
            n_Body_y[278] = c_Body_y[278];
            n_Body_x[279] = c_Body_x[279];
            n_Body_y[279] = c_Body_y[279];
            n_Body_x[280] = c_Body_x[280];
            n_Body_y[280] = c_Body_y[280];
            n_Body_x[281] = c_Body_x[281];
            n_Body_y[281] = c_Body_y[281];
            n_Body_x[282] = c_Body_x[282];
            n_Body_y[282] = c_Body_y[282];
            n_Body_x[283] = c_Body_x[283];
            n_Body_y[283] = c_Body_y[283];
            n_Body_x[284] = c_Body_x[284];
            n_Body_y[284] = c_Body_y[284];
            n_Body_x[285] = c_Body_x[285];
            n_Body_y[285] = c_Body_y[285];
            n_Body_x[286] = c_Body_x[286];
            n_Body_y[286] = c_Body_y[286];
            n_Body_x[287] = c_Body_x[287];
            n_Body_y[287] = c_Body_y[287];
            n_Body_x[288] = c_Body_x[288];
            n_Body_y[288] = c_Body_y[288];
            n_Body_x[289] = c_Body_x[289];
            n_Body_y[289] = c_Body_y[289];
            n_Body_x[290] = c_Body_x[290];
            n_Body_y[290] = c_Body_y[290];
            n_Body_x[291] = c_Body_x[291];
            n_Body_y[291] = c_Body_y[291];
            n_Body_x[292] = c_Body_x[292];
            n_Body_y[292] = c_Body_y[292];
            n_Body_x[293] = c_Body_x[293];
            n_Body_y[293] = c_Body_y[293];
            n_Body_x[294] = c_Body_x[294];
            n_Body_y[294] = c_Body_y[294];
            n_Body_x[295] = c_Body_x[295];
            n_Body_y[295] = c_Body_y[295];
            n_Body_x[296] = c_Body_x[296];
            n_Body_y[296] = c_Body_y[296];
            n_Body_x[297] = c_Body_x[297];
            n_Body_y[297] = c_Body_y[297];
            n_Body_x[298] = c_Body_x[298];
            n_Body_y[298] = c_Body_y[298];
            n_Body_x[299] = c_Body_x[299];
            n_Body_y[299] = c_Body_y[299];
            n_Body_x[300] = c_Body_x[300];
            n_Body_y[300] = c_Body_y[300];
            n_Body_x[301] = c_Body_x[301];
            n_Body_y[301] = c_Body_y[301];
            n_Body_x[302] = c_Body_x[302];
            n_Body_y[302] = c_Body_y[302];
            n_Body_x[303] = c_Body_x[303];
            n_Body_y[303] = c_Body_y[303];
            n_Body_x[304] = c_Body_x[304];
            n_Body_y[304] = c_Body_y[304];
            n_Body_x[305] = c_Body_x[305];
            n_Body_y[305] = c_Body_y[305];
            n_Body_x[306] = c_Body_x[306];
            n_Body_y[306] = c_Body_y[306];
            n_Body_x[307] = c_Body_x[307];
            n_Body_y[307] = c_Body_y[307];
            n_Body_x[308] = c_Body_x[308];
            n_Body_y[308] = c_Body_y[308];
            n_Body_x[309] = c_Body_x[309];
            n_Body_y[309] = c_Body_y[309];
            n_Body_x[310] = c_Body_x[310];
            n_Body_y[310] = c_Body_y[310];
            n_Body_x[311] = c_Body_x[311];
            n_Body_y[311] = c_Body_y[311];
            n_Body_x[312] = c_Body_x[312];
            n_Body_y[312] = c_Body_y[312];
            n_Body_x[313] = c_Body_x[313];
            n_Body_y[313] = c_Body_y[313];
            n_Body_x[314] = c_Body_x[314];
            n_Body_y[314] = c_Body_y[314];
            n_Body_x[315] = c_Body_x[315];
            n_Body_y[315] = c_Body_y[315];
            n_Body_x[316] = c_Body_x[316];
            n_Body_y[316] = c_Body_y[316];
            n_Body_x[317] = c_Body_x[317];
            n_Body_y[317] = c_Body_y[317];
            n_Body_x[318] = c_Body_x[318];
            n_Body_y[318] = c_Body_y[318];
            n_Body_x[319] = c_Body_x[319];
            n_Body_y[319] = c_Body_y[319];
            n_Body_x[320] = c_Body_x[320];
            n_Body_y[320] = c_Body_y[320];
            n_Body_x[321] = c_Body_x[321];
            n_Body_y[321] = c_Body_y[321];
            n_Body_x[322] = c_Body_x[322];
            n_Body_y[322] = c_Body_y[322];
            n_Body_x[323] = c_Body_x[323];
            n_Body_y[323] = c_Body_y[323];
            n_Body_x[324] = c_Body_x[324];
            n_Body_y[324] = c_Body_y[324];
            n_Body_x[325] = c_Body_x[325];
            n_Body_y[325] = c_Body_y[325];
            n_Body_x[326] = c_Body_x[326];
            n_Body_y[326] = c_Body_y[326];
            n_Body_x[327] = c_Body_x[327];
            n_Body_y[327] = c_Body_y[327];
            n_Body_x[328] = c_Body_x[328];
            n_Body_y[328] = c_Body_y[328];
            n_Body_x[329] = c_Body_x[329];
            n_Body_y[329] = c_Body_y[329];
            n_Body_x[330] = c_Body_x[330];
            n_Body_y[330] = c_Body_y[330];
            n_Body_x[331] = c_Body_x[331];
            n_Body_y[331] = c_Body_y[331];
            n_Body_x[332] = c_Body_x[332];
            n_Body_y[332] = c_Body_y[332];
            n_Body_x[333] = c_Body_x[333];
            n_Body_y[333] = c_Body_y[333];
            n_Body_x[334] = c_Body_x[334];
            n_Body_y[334] = c_Body_y[334];
            n_Body_x[335] = c_Body_x[335];
            n_Body_y[335] = c_Body_y[335];
            n_Body_x[336] = c_Body_x[336];
            n_Body_y[336] = c_Body_y[336];
            n_Body_x[337] = c_Body_x[337];
            n_Body_y[337] = c_Body_y[337];
            n_Body_x[338] = c_Body_x[338];
            n_Body_y[338] = c_Body_y[338];
            n_Body_x[339] = c_Body_x[339];
            n_Body_y[339] = c_Body_y[339];
            n_Body_x[340] = c_Body_x[340];
            n_Body_y[340] = c_Body_y[340];
            n_Body_x[341] = c_Body_x[341];
            n_Body_y[341] = c_Body_y[341];
            n_Body_x[342] = c_Body_x[342];
            n_Body_y[342] = c_Body_y[342];
            n_Body_x[343] = c_Body_x[343];
            n_Body_y[343] = c_Body_y[343];
            n_Body_x[344] = c_Body_x[344];
            n_Body_y[344] = c_Body_y[344];
            n_Body_x[345] = c_Body_x[345];
            n_Body_y[345] = c_Body_y[345];
            n_Body_x[346] = c_Body_x[346];
            n_Body_y[346] = c_Body_y[346];
            n_Body_x[347] = c_Body_x[347];
            n_Body_y[347] = c_Body_y[347];
            n_Body_x[348] = c_Body_x[348];
            n_Body_y[348] = c_Body_y[348];
            n_Body_x[349] = c_Body_x[349];
            n_Body_y[349] = c_Body_y[349];
            n_Body_x[350] = c_Body_x[350];
            n_Body_y[350] = c_Body_y[350];
            n_Body_x[351] = c_Body_x[351];
            n_Body_y[351] = c_Body_y[351];
            n_Body_x[352] = c_Body_x[352];
            n_Body_y[352] = c_Body_y[352];
            n_Body_x[353] = c_Body_x[353];
            n_Body_y[353] = c_Body_y[353];
            n_Body_x[354] = c_Body_x[354];
            n_Body_y[354] = c_Body_y[354];
            n_Body_x[355] = c_Body_x[355];
            n_Body_y[355] = c_Body_y[355];
            n_Body_x[356] = c_Body_x[356];
            n_Body_y[356] = c_Body_y[356];
            n_Body_x[357] = c_Body_x[357];
            n_Body_y[357] = c_Body_y[357];
            n_Body_x[358] = c_Body_x[358];
            n_Body_y[358] = c_Body_y[358];
            n_Body_x[359] = c_Body_x[359];
            n_Body_y[359] = c_Body_y[359];
            n_Body_x[360] = c_Body_x[360];
            n_Body_y[360] = c_Body_y[360];
            n_Body_x[361] = c_Body_x[361];
            n_Body_y[361] = c_Body_y[361];
            n_Body_x[362] = c_Body_x[362];
            n_Body_y[362] = c_Body_y[362];
            n_Body_x[363] = c_Body_x[363];
            n_Body_y[363] = c_Body_y[363];
            n_Body_x[364] = c_Body_x[364];
            n_Body_y[364] = c_Body_y[364];
            n_Body_x[365] = c_Body_x[365];
            n_Body_y[365] = c_Body_y[365];
            n_Body_x[366] = c_Body_x[366];
            n_Body_y[366] = c_Body_y[366];
            n_Body_x[367] = c_Body_x[367];
            n_Body_y[367] = c_Body_y[367];
            n_Body_x[368] = c_Body_x[368];
            n_Body_y[368] = c_Body_y[368];
            n_Body_x[369] = c_Body_x[369];
            n_Body_y[369] = c_Body_y[369];
            n_Body_x[370] = c_Body_x[370];
            n_Body_y[370] = c_Body_y[370];
            n_Body_x[371] = c_Body_x[371];
            n_Body_y[371] = c_Body_y[371];
            n_Body_x[372] = c_Body_x[372];
            n_Body_y[372] = c_Body_y[372];
            n_Body_x[373] = c_Body_x[373];
            n_Body_y[373] = c_Body_y[373];
            n_Body_x[374] = c_Body_x[374];
            n_Body_y[374] = c_Body_y[374];
            n_Body_x[375] = c_Body_x[375];
            n_Body_y[375] = c_Body_y[375];
            n_Body_x[376] = c_Body_x[376];
            n_Body_y[376] = c_Body_y[376];
            n_Body_x[377] = c_Body_x[377];
            n_Body_y[377] = c_Body_y[377];
            n_Body_x[378] = c_Body_x[378];
            n_Body_y[378] = c_Body_y[378];
            n_Body_x[379] = c_Body_x[379];
            n_Body_y[379] = c_Body_y[379];
            n_Body_x[380] = c_Body_x[380];
            n_Body_y[380] = c_Body_y[380];
            n_Body_x[381] = c_Body_x[381];
            n_Body_y[381] = c_Body_y[381];
            n_Body_x[382] = c_Body_x[382];
            n_Body_y[382] = c_Body_y[382];
            n_Body_x[383] = c_Body_x[383];
            n_Body_y[383] = c_Body_y[383];
            n_Body_x[384] = c_Body_x[384];
            n_Body_y[384] = c_Body_y[384];
            n_Body_x[385] = c_Body_x[385];
            n_Body_y[385] = c_Body_y[385];
            n_Body_x[386] = c_Body_x[386];
            n_Body_y[386] = c_Body_y[386];
            n_Body_x[387] = c_Body_x[387];
            n_Body_y[387] = c_Body_y[387];
            n_Body_x[388] = c_Body_x[388];
            n_Body_y[388] = c_Body_y[388];
            n_Body_x[389] = c_Body_x[389];
            n_Body_y[389] = c_Body_y[389];
            n_Body_x[390] = c_Body_x[390];
            n_Body_y[390] = c_Body_y[390];
            n_Body_x[391] = c_Body_x[391];
            n_Body_y[391] = c_Body_y[391];
            n_Body_x[392] = c_Body_x[392];
            n_Body_y[392] = c_Body_y[392];
            n_Body_x[393] = c_Body_x[393];
            n_Body_y[393] = c_Body_y[393];
            n_Body_x[394] = c_Body_x[394];
            n_Body_y[394] = c_Body_y[394];
            n_Body_x[395] = c_Body_x[395];
            n_Body_y[395] = c_Body_y[395];
            n_Body_x[396] = c_Body_x[396];
            n_Body_y[396] = c_Body_y[396];
            n_Body_x[397] = c_Body_x[397];
            n_Body_y[397] = c_Body_y[397];
            n_Body_x[398] = c_Body_x[398];
            n_Body_y[398] = c_Body_y[398];
            n_Body_x[399] = c_Body_x[399];
            n_Body_y[399] = c_Body_y[399];
            n_Body_x[400] = c_Body_x[400];
            n_Body_y[400] = c_Body_y[400];
            n_Body_x[401] = c_Body_x[401];
            n_Body_y[401] = c_Body_y[401];
            n_Body_x[402] = c_Body_x[402];
            n_Body_y[402] = c_Body_y[402];
            n_Body_x[403] = c_Body_x[403];
            n_Body_y[403] = c_Body_y[403];
            n_Body_x[404] = c_Body_x[404];
            n_Body_y[404] = c_Body_y[404];
            n_Body_x[405] = c_Body_x[405];
            n_Body_y[405] = c_Body_y[405];
            n_Body_x[406] = c_Body_x[406];
            n_Body_y[406] = c_Body_y[406];
            n_Body_x[407] = c_Body_x[407];
            n_Body_y[407] = c_Body_y[407];
            n_Body_x[408] = c_Body_x[408];
            n_Body_y[408] = c_Body_y[408];
            n_Body_x[409] = c_Body_x[409];
            n_Body_y[409] = c_Body_y[409];
            n_Body_x[410] = c_Body_x[410];
            n_Body_y[410] = c_Body_y[410];
            n_Body_x[411] = c_Body_x[411];
            n_Body_y[411] = c_Body_y[411];
            n_Body_x[412] = c_Body_x[412];
            n_Body_y[412] = c_Body_y[412];
            n_Body_x[413] = c_Body_x[413];
            n_Body_y[413] = c_Body_y[413];
            n_Body_x[414] = c_Body_x[414];
            n_Body_y[414] = c_Body_y[414];
            n_Body_x[415] = c_Body_x[415];
            n_Body_y[415] = c_Body_y[415];
            n_Body_x[416] = c_Body_x[416];
            n_Body_y[416] = c_Body_y[416];
            n_Body_x[417] = c_Body_x[417];
            n_Body_y[417] = c_Body_y[417];
            n_Body_x[418] = c_Body_x[418];
            n_Body_y[418] = c_Body_y[418];
            n_Body_x[419] = c_Body_x[419];
            n_Body_y[419] = c_Body_y[419];
            n_Body_x[420] = c_Body_x[420];
            n_Body_y[420] = c_Body_y[420];
            n_Body_x[421] = c_Body_x[421];
            n_Body_y[421] = c_Body_y[421];
            n_Body_x[422] = c_Body_x[422];
            n_Body_y[422] = c_Body_y[422];
            n_Body_x[423] = c_Body_x[423];
            n_Body_y[423] = c_Body_y[423];
            n_Body_x[424] = c_Body_x[424];
            n_Body_y[424] = c_Body_y[424];
            n_Body_x[425] = c_Body_x[425];
            n_Body_y[425] = c_Body_y[425];
            n_Body_x[426] = c_Body_x[426];
            n_Body_y[426] = c_Body_y[426];
            n_Body_x[427] = c_Body_x[427];
            n_Body_y[427] = c_Body_y[427];
            n_Body_x[428] = c_Body_x[428];
            n_Body_y[428] = c_Body_y[428];
            n_Body_x[429] = c_Body_x[429];
            n_Body_y[429] = c_Body_y[429];
            n_Body_x[430] = c_Body_x[430];
            n_Body_y[430] = c_Body_y[430];
            n_Body_x[431] = c_Body_x[431];
            n_Body_y[431] = c_Body_y[431];
            n_Body_x[432] = c_Body_x[432];
            n_Body_y[432] = c_Body_y[432];
            n_Body_x[433] = c_Body_x[433];
            n_Body_y[433] = c_Body_y[433];
            n_Body_x[434] = c_Body_x[434];
            n_Body_y[434] = c_Body_y[434];
            n_Body_x[435] = c_Body_x[435];
            n_Body_y[435] = c_Body_y[435];
            n_Body_x[436] = c_Body_x[436];
            n_Body_y[436] = c_Body_y[436];
            n_Body_x[437] = c_Body_x[437];
            n_Body_y[437] = c_Body_y[437];
            n_Body_x[438] = c_Body_x[438];
            n_Body_y[438] = c_Body_y[438];
            n_Body_x[439] = c_Body_x[439];
            n_Body_y[439] = c_Body_y[439];
            n_Body_x[440] = c_Body_x[440];
            n_Body_y[440] = c_Body_y[440];
            n_Body_x[441] = c_Body_x[441];
            n_Body_y[441] = c_Body_y[441];
            n_Body_x[442] = c_Body_x[442];
            n_Body_y[442] = c_Body_y[442];
            n_Body_x[443] = c_Body_x[443];
            n_Body_y[443] = c_Body_y[443];
            n_Body_x[444] = c_Body_x[444];
            n_Body_y[444] = c_Body_y[444];
            n_Body_x[445] = c_Body_x[445];
            n_Body_y[445] = c_Body_y[445];
            n_Body_x[446] = c_Body_x[446];
            n_Body_y[446] = c_Body_y[446];
            n_Body_x[447] = c_Body_x[447];
            n_Body_y[447] = c_Body_y[447];
            n_Body_x[448] = c_Body_x[448];
            n_Body_y[448] = c_Body_y[448];
            n_Body_x[449] = c_Body_x[449];
            n_Body_y[449] = c_Body_y[449];
            n_Body_x[450] = c_Body_x[450];
            n_Body_y[450] = c_Body_y[450];
            n_Body_x[451] = c_Body_x[451];
            n_Body_y[451] = c_Body_y[451];
            n_Body_x[452] = c_Body_x[452];
            n_Body_y[452] = c_Body_y[452];
            n_Body_x[453] = c_Body_x[453];
            n_Body_y[453] = c_Body_y[453];
            n_Body_x[454] = c_Body_x[454];
            n_Body_y[454] = c_Body_y[454];
            n_Body_x[455] = c_Body_x[455];
            n_Body_y[455] = c_Body_y[455];
            n_Body_x[456] = c_Body_x[456];
            n_Body_y[456] = c_Body_y[456];
            n_Body_x[457] = c_Body_x[457];
            n_Body_y[457] = c_Body_y[457];
            n_Body_x[458] = c_Body_x[458];
            n_Body_y[458] = c_Body_y[458];
            n_Body_x[459] = c_Body_x[459];
            n_Body_y[459] = c_Body_y[459];
            n_Body_x[460] = c_Body_x[460];
            n_Body_y[460] = c_Body_y[460];
            n_Body_x[461] = c_Body_x[461];
            n_Body_y[461] = c_Body_y[461];
            n_Body_x[462] = c_Body_x[462];
            n_Body_y[462] = c_Body_y[462];
            n_Body_x[463] = c_Body_x[463];
            n_Body_y[463] = c_Body_y[463];
            n_Body_x[464] = c_Body_x[464];
            n_Body_y[464] = c_Body_y[464];
            n_Body_x[465] = c_Body_x[465];
            n_Body_y[465] = c_Body_y[465];
            n_Body_x[466] = c_Body_x[466];
            n_Body_y[466] = c_Body_y[466];
            n_Body_x[467] = c_Body_x[467];
            n_Body_y[467] = c_Body_y[467];
            n_Body_x[468] = c_Body_x[468];
            n_Body_y[468] = c_Body_y[468];
            n_Body_x[469] = c_Body_x[469];
            n_Body_y[469] = c_Body_y[469];
            n_Body_x[470] = c_Body_x[470];
            n_Body_y[470] = c_Body_y[470];
            n_Body_x[471] = c_Body_x[471];
            n_Body_y[471] = c_Body_y[471];
            n_Body_x[472] = c_Body_x[472];
            n_Body_y[472] = c_Body_y[472];
            n_Body_x[473] = c_Body_x[473];
            n_Body_y[473] = c_Body_y[473];
            n_Body_x[474] = c_Body_x[474];
            n_Body_y[474] = c_Body_y[474];
            n_Body_x[475] = c_Body_x[475];
            n_Body_y[475] = c_Body_y[475];
            n_Body_x[476] = c_Body_x[476];
            n_Body_y[476] = c_Body_y[476];
            n_Body_x[477] = c_Body_x[477];
            n_Body_y[477] = c_Body_y[477];
            n_Body_x[478] = c_Body_x[478];
            n_Body_y[478] = c_Body_y[478];
            n_Body_x[479] = c_Body_x[479];
            n_Body_y[479] = c_Body_y[479];
            n_Body_x[480] = c_Body_x[480];
            n_Body_y[480] = c_Body_y[480];
            n_Body_x[481] = c_Body_x[481];
            n_Body_y[481] = c_Body_y[481];
            n_Body_x[482] = c_Body_x[482];
            n_Body_y[482] = c_Body_y[482];
            n_Body_x[483] = c_Body_x[483];
            n_Body_y[483] = c_Body_y[483];
            n_Body_x[484] = c_Body_x[484];
            n_Body_y[484] = c_Body_y[484];
            n_Body_x[485] = c_Body_x[485];
            n_Body_y[485] = c_Body_y[485];
            n_Body_x[486] = c_Body_x[486];
            n_Body_y[486] = c_Body_y[486];
            n_Body_x[487] = c_Body_x[487];
            n_Body_y[487] = c_Body_y[487];
            n_Body_x[488] = c_Body_x[488];
            n_Body_y[488] = c_Body_y[488];
            n_Body_x[489] = c_Body_x[489];
            n_Body_y[489] = c_Body_y[489];
            n_Body_x[490] = c_Body_x[490];
            n_Body_y[490] = c_Body_y[490];
            n_Body_x[491] = c_Body_x[491];
            n_Body_y[491] = c_Body_y[491];
            n_Body_x[492] = c_Body_x[492];
            n_Body_y[492] = c_Body_y[492];
            n_Body_x[493] = c_Body_x[493];
            n_Body_y[493] = c_Body_y[493];
            n_Body_x[494] = c_Body_x[494];
            n_Body_y[494] = c_Body_y[494];
            n_Body_x[495] = c_Body_x[495];
            n_Body_y[495] = c_Body_y[495];
            n_Body_x[496] = c_Body_x[496];
            n_Body_y[496] = c_Body_y[496];
            n_Body_x[497] = c_Body_x[497];
            n_Body_y[497] = c_Body_y[497];
            n_Body_x[498] = c_Body_x[498];
            n_Body_y[498] = c_Body_y[498];
            n_Body_x[499] = c_Body_x[499];
            n_Body_y[499] = c_Body_y[499];
            n_Body_x[500] = c_Body_x[500];
            n_Body_y[500] = c_Body_y[500];
            n_Body_x[501] = c_Body_x[501];
            n_Body_y[501] = c_Body_y[501];
            n_Body_x[502] = c_Body_x[502];
            n_Body_y[502] = c_Body_y[502];
            n_Body_x[503] = c_Body_x[503];
            n_Body_y[503] = c_Body_y[503];
            n_Body_x[504] = c_Body_x[504];
            n_Body_y[504] = c_Body_y[504];
            n_Body_x[505] = c_Body_x[505];
            n_Body_y[505] = c_Body_y[505];
            n_Body_x[506] = c_Body_x[506];
            n_Body_y[506] = c_Body_y[506];
            n_Body_x[507] = c_Body_x[507];
            n_Body_y[507] = c_Body_y[507];
            n_Body_x[508] = c_Body_x[508];
            n_Body_y[508] = c_Body_y[508];
            n_Body_x[509] = c_Body_x[509];
            n_Body_y[509] = c_Body_y[509];
            n_Body_x[510] = c_Body_x[510];
            n_Body_y[510] = c_Body_y[510];
            n_Body_x[511] = c_Body_x[511];
            n_Body_y[511] = c_Body_y[511];
            n_Body_x[512] = c_Body_x[512];
            n_Body_y[512] = c_Body_y[512];
            n_Body_x[513] = c_Body_x[513];
            n_Body_y[513] = c_Body_y[513];
            n_Body_x[514] = c_Body_x[514];
            n_Body_y[514] = c_Body_y[514];
            n_Body_x[515] = c_Body_x[515];
            n_Body_y[515] = c_Body_y[515];
            n_Body_x[516] = c_Body_x[516];
            n_Body_y[516] = c_Body_y[516];
            n_Body_x[517] = c_Body_x[517];
            n_Body_y[517] = c_Body_y[517];
            n_Body_x[518] = c_Body_x[518];
            n_Body_y[518] = c_Body_y[518];
            n_Body_x[519] = c_Body_x[519];
            n_Body_y[519] = c_Body_y[519];
            n_Body_x[520] = c_Body_x[520];
            n_Body_y[520] = c_Body_y[520];
            n_Body_x[521] = c_Body_x[521];
            n_Body_y[521] = c_Body_y[521];
            n_Body_x[522] = c_Body_x[522];
            n_Body_y[522] = c_Body_y[522];
            n_Body_x[523] = c_Body_x[523];
            n_Body_y[523] = c_Body_y[523];
            n_Body_x[524] = c_Body_x[524];
            n_Body_y[524] = c_Body_y[524];
            n_Body_x[525] = c_Body_x[525];
            n_Body_y[525] = c_Body_y[525];
            n_Body_x[526] = c_Body_x[526];
            n_Body_y[526] = c_Body_y[526];
            n_Body_x[527] = c_Body_x[527];
            n_Body_y[527] = c_Body_y[527];
            n_Body_x[528] = c_Body_x[528];
            n_Body_y[528] = c_Body_y[528];
            n_Body_x[529] = c_Body_x[529];
            n_Body_y[529] = c_Body_y[529];
            n_Body_x[530] = c_Body_x[530];
            n_Body_y[530] = c_Body_y[530];
            n_Body_x[531] = c_Body_x[531];
            n_Body_y[531] = c_Body_y[531];
            n_Body_x[532] = c_Body_x[532];
            n_Body_y[532] = c_Body_y[532];
            n_Body_x[533] = c_Body_x[533];
            n_Body_y[533] = c_Body_y[533];
            n_Body_x[534] = c_Body_x[534];
            n_Body_y[534] = c_Body_y[534];
            n_Body_x[535] = c_Body_x[535];
            n_Body_y[535] = c_Body_y[535];
            n_Body_x[536] = c_Body_x[536];
            n_Body_y[536] = c_Body_y[536];
            n_Body_x[537] = c_Body_x[537];
            n_Body_y[537] = c_Body_y[537];
            n_Body_x[538] = c_Body_x[538];
            n_Body_y[538] = c_Body_y[538];
            n_Body_x[539] = c_Body_x[539];
            n_Body_y[539] = c_Body_y[539];
            n_Body_x[540] = c_Body_x[540];
            n_Body_y[540] = c_Body_y[540];
            n_Body_x[541] = c_Body_x[541];
            n_Body_y[541] = c_Body_y[541];
            n_Body_x[542] = c_Body_x[542];
            n_Body_y[542] = c_Body_y[542];
            n_Body_x[543] = c_Body_x[543];
            n_Body_y[543] = c_Body_y[543];
            n_Body_x[544] = c_Body_x[544];
            n_Body_y[544] = c_Body_y[544];
            n_Body_x[545] = c_Body_x[545];
            n_Body_y[545] = c_Body_y[545];
            n_Body_x[546] = c_Body_x[546];
            n_Body_y[546] = c_Body_y[546];
            n_Body_x[547] = c_Body_x[547];
            n_Body_y[547] = c_Body_y[547];
            n_Body_x[548] = c_Body_x[548];
            n_Body_y[548] = c_Body_y[548];
            n_Body_x[549] = c_Body_x[549];
            n_Body_y[549] = c_Body_y[549];
            n_Body_x[550] = c_Body_x[550];
            n_Body_y[550] = c_Body_y[550];
            n_Body_x[551] = c_Body_x[551];
            n_Body_y[551] = c_Body_y[551];
            n_Body_x[552] = c_Body_x[552];
            n_Body_y[552] = c_Body_y[552];
            n_Body_x[553] = c_Body_x[553];
            n_Body_y[553] = c_Body_y[553];
            n_Body_x[554] = c_Body_x[554];
            n_Body_y[554] = c_Body_y[554];
            n_Body_x[555] = c_Body_x[555];
            n_Body_y[555] = c_Body_y[555];
            n_Body_x[556] = c_Body_x[556];
            n_Body_y[556] = c_Body_y[556];
            n_Body_x[557] = c_Body_x[557];
            n_Body_y[557] = c_Body_y[557];
            n_Body_x[558] = c_Body_x[558];
            n_Body_y[558] = c_Body_y[558];
            n_Body_x[559] = c_Body_x[559];
            n_Body_y[559] = c_Body_y[559];
            n_Body_x[560] = c_Body_x[560];
            n_Body_y[560] = c_Body_y[560];
            n_Body_x[561] = c_Body_x[561];
            n_Body_y[561] = c_Body_y[561];
            n_Body_x[562] = c_Body_x[562];
            n_Body_y[562] = c_Body_y[562];
            n_Body_x[563] = c_Body_x[563];
            n_Body_y[563] = c_Body_y[563];
            n_Body_x[564] = c_Body_x[564];
            n_Body_y[564] = c_Body_y[564];
            n_Body_x[565] = c_Body_x[565];
            n_Body_y[565] = c_Body_y[565];
            n_Body_x[566] = c_Body_x[566];
            n_Body_y[566] = c_Body_y[566];
            n_Body_x[567] = c_Body_x[567];
            n_Body_y[567] = c_Body_y[567];
            n_Body_x[568] = c_Body_x[568];
            n_Body_y[568] = c_Body_y[568];
            n_Body_x[569] = c_Body_x[569];
            n_Body_y[569] = c_Body_y[569];
            n_Body_x[570] = c_Body_x[570];
            n_Body_y[570] = c_Body_y[570];
            n_Body_x[571] = c_Body_x[571];
            n_Body_y[571] = c_Body_y[571];
            n_Body_x[572] = c_Body_x[572];
            n_Body_y[572] = c_Body_y[572];
            n_Body_x[573] = c_Body_x[573];
            n_Body_y[573] = c_Body_y[573];
            n_Body_x[574] = c_Body_x[574];
            n_Body_y[574] = c_Body_y[574];
            n_Body_x[575] = c_Body_x[575];
            n_Body_y[575] = c_Body_y[575];
            n_Body_x[576] = c_Body_x[576];
            n_Body_y[576] = c_Body_y[576];
            n_Body_x[577] = c_Body_x[577];
            n_Body_y[577] = c_Body_y[577];
            n_Body_x[578] = c_Body_x[578];
            n_Body_y[578] = c_Body_y[578];
            n_Body_x[579] = c_Body_x[579];
            n_Body_y[579] = c_Body_y[579];
            n_Body_x[580] = c_Body_x[580];
            n_Body_y[580] = c_Body_y[580];
            n_Body_x[581] = c_Body_x[581];
            n_Body_y[581] = c_Body_y[581];
            n_Body_x[582] = c_Body_x[582];
            n_Body_y[582] = c_Body_y[582];
            n_Body_x[583] = c_Body_x[583];
            n_Body_y[583] = c_Body_y[583];
            n_Body_x[584] = c_Body_x[584];
            n_Body_y[584] = c_Body_y[584];
            n_Body_x[585] = c_Body_x[585];
            n_Body_y[585] = c_Body_y[585];
            n_Body_x[586] = c_Body_x[586];
            n_Body_y[586] = c_Body_y[586];
            n_Body_x[587] = c_Body_x[587];
            n_Body_y[587] = c_Body_y[587];
            n_Body_x[588] = c_Body_x[588];
            n_Body_y[588] = c_Body_y[588];
            n_Body_x[589] = c_Body_x[589];
            n_Body_y[589] = c_Body_y[589];
            n_Body_x[590] = c_Body_x[590];
            n_Body_y[590] = c_Body_y[590];
            n_Body_x[591] = c_Body_x[591];
            n_Body_y[591] = c_Body_y[591];
            n_Body_x[592] = c_Body_x[592];
            n_Body_y[592] = c_Body_y[592];
            n_Body_x[593] = c_Body_x[593];
            n_Body_y[593] = c_Body_y[593];
            n_Body_x[594] = c_Body_x[594];
            n_Body_y[594] = c_Body_y[594];
            n_Body_x[595] = c_Body_x[595];
            n_Body_y[595] = c_Body_y[595];
            n_Body_x[596] = c_Body_x[596];
            n_Body_y[596] = c_Body_y[596];
            n_Body_x[597] = c_Body_x[597];
            n_Body_y[597] = c_Body_y[597];
            n_Body_x[598] = c_Body_x[598];
            n_Body_y[598] = c_Body_y[598];
            n_Body_x[599] = c_Body_x[599];
            n_Body_y[599] = c_Body_y[599];
            n_Body_x[600] = c_Body_x[600];
            n_Body_y[600] = c_Body_y[600];
            n_Body_x[601] = c_Body_x[601];
            n_Body_y[601] = c_Body_y[601];
            n_Body_x[602] = c_Body_x[602];
            n_Body_y[602] = c_Body_y[602];
            n_Body_x[603] = c_Body_x[603];
            n_Body_y[603] = c_Body_y[603];
            n_Body_x[604] = c_Body_x[604];
            n_Body_y[604] = c_Body_y[604];
            n_Body_x[605] = c_Body_x[605];
            n_Body_y[605] = c_Body_y[605];
            n_Body_x[606] = c_Body_x[606];
            n_Body_y[606] = c_Body_y[606];
            n_Body_x[607] = c_Body_x[607];
            n_Body_y[607] = c_Body_y[607];
            n_Body_x[608] = c_Body_x[608];
            n_Body_y[608] = c_Body_y[608];
            n_Body_x[609] = c_Body_x[609];
            n_Body_y[609] = c_Body_y[609];
            n_Body_x[610] = c_Body_x[610];
            n_Body_y[610] = c_Body_y[610];
            n_Body_x[611] = c_Body_x[611];
            n_Body_y[611] = c_Body_y[611];
            n_Body_x[612] = c_Body_x[612];
            n_Body_y[612] = c_Body_y[612];
            n_Body_x[613] = c_Body_x[613];
            n_Body_y[613] = c_Body_y[613];
            n_Body_x[614] = c_Body_x[614];
            n_Body_y[614] = c_Body_y[614];
            n_Body_x[615] = c_Body_x[615];
            n_Body_y[615] = c_Body_y[615];
            n_Body_x[616] = c_Body_x[616];
            n_Body_y[616] = c_Body_y[616];
            n_Body_x[617] = c_Body_x[617];
            n_Body_y[617] = c_Body_y[617];
            n_Body_x[618] = c_Body_x[618];
            n_Body_y[618] = c_Body_y[618];
            n_Body_x[619] = c_Body_x[619];
            n_Body_y[619] = c_Body_y[619];
            n_Body_x[620] = c_Body_x[620];
            n_Body_y[620] = c_Body_y[620];
            n_Body_x[621] = c_Body_x[621];
            n_Body_y[621] = c_Body_y[621];
            n_Body_x[622] = c_Body_x[622];
            n_Body_y[622] = c_Body_y[622];
            n_Body_x[623] = c_Body_x[623];
            n_Body_y[623] = c_Body_y[623];
            n_Body_x[624] = c_Body_x[624];
            n_Body_y[624] = c_Body_y[624];
            n_Body_x[625] = c_Body_x[625];
            n_Body_y[625] = c_Body_y[625];
            n_Body_x[626] = c_Body_x[626];
            n_Body_y[626] = c_Body_y[626];
            n_Body_x[627] = c_Body_x[627];
            n_Body_y[627] = c_Body_y[627];
            n_Body_x[628] = c_Body_x[628];
            n_Body_y[628] = c_Body_y[628];
            n_Body_x[629] = c_Body_x[629];
            n_Body_y[629] = c_Body_y[629];
            n_Body_x[630] = c_Body_x[630];
            n_Body_y[630] = c_Body_y[630];
            n_Body_x[631] = c_Body_x[631];
            n_Body_y[631] = c_Body_y[631];
            n_Body_x[632] = c_Body_x[632];
            n_Body_y[632] = c_Body_y[632];
            n_Body_x[633] = c_Body_x[633];
            n_Body_y[633] = c_Body_y[633];
            n_Body_x[634] = c_Body_x[634];
            n_Body_y[634] = c_Body_y[634];
            n_Body_x[635] = c_Body_x[635];
            n_Body_y[635] = c_Body_y[635];
            n_Body_x[636] = c_Body_x[636];
            n_Body_y[636] = c_Body_y[636];
            n_Body_x[637] = c_Body_x[637];
            n_Body_y[637] = c_Body_y[637];
            n_Body_x[638] = c_Body_x[638];
            n_Body_y[638] = c_Body_y[638];
            n_Body_x[639] = c_Body_x[639];
            n_Body_y[639] = c_Body_y[639];
            n_Body_x[640] = c_Body_x[640];
            n_Body_y[640] = c_Body_y[640];
            n_Body_x[641] = c_Body_x[641];
            n_Body_y[641] = c_Body_y[641];
            n_Body_x[642] = c_Body_x[642];
            n_Body_y[642] = c_Body_y[642];
            n_Body_x[643] = c_Body_x[643];
            n_Body_y[643] = c_Body_y[643];
            n_Body_x[644] = c_Body_x[644];
            n_Body_y[644] = c_Body_y[644];
            n_Body_x[645] = c_Body_x[645];
            n_Body_y[645] = c_Body_y[645];
            n_Body_x[646] = c_Body_x[646];
            n_Body_y[646] = c_Body_y[646];
            n_Body_x[647] = c_Body_x[647];
            n_Body_y[647] = c_Body_y[647];
            n_Body_x[648] = c_Body_x[648];
            n_Body_y[648] = c_Body_y[648];
            n_Body_x[649] = c_Body_x[649];
            n_Body_y[649] = c_Body_y[649];
            n_Body_x[650] = c_Body_x[650];
            n_Body_y[650] = c_Body_y[650];
            n_Body_x[651] = c_Body_x[651];
            n_Body_y[651] = c_Body_y[651];
            n_Body_x[652] = c_Body_x[652];
            n_Body_y[652] = c_Body_y[652];
            n_Body_x[653] = c_Body_x[653];
            n_Body_y[653] = c_Body_y[653];
            n_Body_x[654] = c_Body_x[654];
            n_Body_y[654] = c_Body_y[654];
            n_Body_x[655] = c_Body_x[655];
            n_Body_y[655] = c_Body_y[655];
            n_Body_x[656] = c_Body_x[656];
            n_Body_y[656] = c_Body_y[656];
            n_Body_x[657] = c_Body_x[657];
            n_Body_y[657] = c_Body_y[657];
            n_Body_x[658] = c_Body_x[658];
            n_Body_y[658] = c_Body_y[658];
            n_Body_x[659] = c_Body_x[659];
            n_Body_y[659] = c_Body_y[659];
            n_Body_x[660] = c_Body_x[660];
            n_Body_y[660] = c_Body_y[660];
            n_Body_x[661] = c_Body_x[661];
            n_Body_y[661] = c_Body_y[661];
            n_Body_x[662] = c_Body_x[662];
            n_Body_y[662] = c_Body_y[662];
            n_Body_x[663] = c_Body_x[663];
            n_Body_y[663] = c_Body_y[663];
            n_Body_x[664] = c_Body_x[664];
            n_Body_y[664] = c_Body_y[664];
            n_Body_x[665] = c_Body_x[665];
            n_Body_y[665] = c_Body_y[665];
            n_Body_x[666] = c_Body_x[666];
            n_Body_y[666] = c_Body_y[666];
            n_Body_x[667] = c_Body_x[667];
            n_Body_y[667] = c_Body_y[667];
            n_Body_x[668] = c_Body_x[668];
            n_Body_y[668] = c_Body_y[668];
            n_Body_x[669] = c_Body_x[669];
            n_Body_y[669] = c_Body_y[669];
            n_Body_x[670] = c_Body_x[670];
            n_Body_y[670] = c_Body_y[670];
            n_Body_x[671] = c_Body_x[671];
            n_Body_y[671] = c_Body_y[671];
            n_Body_x[672] = c_Body_x[672];
            n_Body_y[672] = c_Body_y[672];
            n_Body_x[673] = c_Body_x[673];
            n_Body_y[673] = c_Body_y[673];
            n_Body_x[674] = c_Body_x[674];
            n_Body_y[674] = c_Body_y[674];
            n_Body_x[675] = c_Body_x[675];
            n_Body_y[675] = c_Body_y[675];
            n_Body_x[676] = c_Body_x[676];
            n_Body_y[676] = c_Body_y[676];
            n_Body_x[677] = c_Body_x[677];
            n_Body_y[677] = c_Body_y[677];
            n_Body_x[678] = c_Body_x[678];
            n_Body_y[678] = c_Body_y[678];
            n_Body_x[679] = c_Body_x[679];
            n_Body_y[679] = c_Body_y[679];
            n_Body_x[680] = c_Body_x[680];
            n_Body_y[680] = c_Body_y[680];
            n_Body_x[681] = c_Body_x[681];
            n_Body_y[681] = c_Body_y[681];
            n_Body_x[682] = c_Body_x[682];
            n_Body_y[682] = c_Body_y[682];
            n_Body_x[683] = c_Body_x[683];
            n_Body_y[683] = c_Body_y[683];
            n_Body_x[684] = c_Body_x[684];
            n_Body_y[684] = c_Body_y[684];
            n_Body_x[685] = c_Body_x[685];
            n_Body_y[685] = c_Body_y[685];
            n_Body_x[686] = c_Body_x[686];
            n_Body_y[686] = c_Body_y[686];
            n_Body_x[687] = c_Body_x[687];
            n_Body_y[687] = c_Body_y[687];
            n_Body_x[688] = c_Body_x[688];
            n_Body_y[688] = c_Body_y[688];
            n_Body_x[689] = c_Body_x[689];
            n_Body_y[689] = c_Body_y[689];
            n_Body_x[690] = c_Body_x[690];
            n_Body_y[690] = c_Body_y[690];
            n_Body_x[691] = c_Body_x[691];
            n_Body_y[691] = c_Body_y[691];
            n_Body_x[692] = c_Body_x[692];
            n_Body_y[692] = c_Body_y[692];
            n_Body_x[693] = c_Body_x[693];
            n_Body_y[693] = c_Body_y[693];
            n_Body_x[694] = c_Body_x[694];
            n_Body_y[694] = c_Body_y[694];
            n_Body_x[695] = c_Body_x[695];
            n_Body_y[695] = c_Body_y[695];
            n_Body_x[696] = c_Body_x[696];
            n_Body_y[696] = c_Body_y[696];
            n_Body_x[697] = c_Body_x[697];
            n_Body_y[697] = c_Body_y[697];
            n_Body_x[698] = c_Body_x[698];
            n_Body_y[698] = c_Body_y[698];
            n_Body_x[699] = c_Body_x[699];
            n_Body_y[699] = c_Body_y[699];
            n_Body_x[700] = c_Body_x[700];
            n_Body_y[700] = c_Body_y[700];
            n_Body_x[701] = c_Body_x[701];
            n_Body_y[701] = c_Body_y[701];
            n_Body_x[702] = c_Body_x[702];
            n_Body_y[702] = c_Body_y[702];
            n_Body_x[703] = c_Body_x[703];
            n_Body_y[703] = c_Body_y[703];
            n_Body_x[704] = c_Body_x[704];
            n_Body_y[704] = c_Body_y[704];
            n_Body_x[705] = c_Body_x[705];
            n_Body_y[705] = c_Body_y[705];
            n_Body_x[706] = c_Body_x[706];
            n_Body_y[706] = c_Body_y[706];
            n_Body_x[707] = c_Body_x[707];
            n_Body_y[707] = c_Body_y[707];
            n_Body_x[708] = c_Body_x[708];
            n_Body_y[708] = c_Body_y[708];
            n_Body_x[709] = c_Body_x[709];
            n_Body_y[709] = c_Body_y[709];
            n_Body_x[710] = c_Body_x[710];
            n_Body_y[710] = c_Body_y[710];
            n_Body_x[711] = c_Body_x[711];
            n_Body_y[711] = c_Body_y[711];
            n_Body_x[712] = c_Body_x[712];
            n_Body_y[712] = c_Body_y[712];
            n_Body_x[713] = c_Body_x[713];
            n_Body_y[713] = c_Body_y[713];
            n_Body_x[714] = c_Body_x[714];
            n_Body_y[714] = c_Body_y[714];
            n_Body_x[715] = c_Body_x[715];
            n_Body_y[715] = c_Body_y[715];
            n_Body_x[716] = c_Body_x[716];
            n_Body_y[716] = c_Body_y[716];
            n_Body_x[717] = c_Body_x[717];
            n_Body_y[717] = c_Body_y[717];
            n_Body_x[718] = c_Body_x[718];
            n_Body_y[718] = c_Body_y[718];
            n_Body_x[719] = c_Body_x[719];
            n_Body_y[719] = c_Body_y[719];
            n_Body_x[720] = c_Body_x[720];
            n_Body_y[720] = c_Body_y[720];
            n_Body_x[721] = c_Body_x[721];
            n_Body_y[721] = c_Body_y[721];
            n_Body_x[722] = c_Body_x[722];
            n_Body_y[722] = c_Body_y[722];
            n_Body_x[723] = c_Body_x[723];
            n_Body_y[723] = c_Body_y[723];
            n_Body_x[724] = c_Body_x[724];
            n_Body_y[724] = c_Body_y[724];
            n_Body_x[725] = c_Body_x[725];
            n_Body_y[725] = c_Body_y[725];
            n_Body_x[726] = c_Body_x[726];
            n_Body_y[726] = c_Body_y[726];
            n_Body_x[727] = c_Body_x[727];
            n_Body_y[727] = c_Body_y[727];
            n_Body_x[728] = c_Body_x[728];
            n_Body_y[728] = c_Body_y[728];
            n_Body_x[729] = c_Body_x[729];
            n_Body_y[729] = c_Body_y[729];
            n_Body_x[730] = c_Body_x[730];
            n_Body_y[730] = c_Body_y[730];
            n_Body_x[731] = c_Body_x[731];
            n_Body_y[731] = c_Body_y[731];
            n_Body_x[732] = c_Body_x[732];
            n_Body_y[732] = c_Body_y[732];
            n_Body_x[733] = c_Body_x[733];
            n_Body_y[733] = c_Body_y[733];
            n_Body_x[734] = c_Body_x[734];
            n_Body_y[734] = c_Body_y[734];
            n_Body_x[735] = c_Body_x[735];
            n_Body_y[735] = c_Body_y[735];
            n_Body_x[736] = c_Body_x[736];
            n_Body_y[736] = c_Body_y[736];
            n_Body_x[737] = c_Body_x[737];
            n_Body_y[737] = c_Body_y[737];
            n_Body_x[738] = c_Body_x[738];
            n_Body_y[738] = c_Body_y[738];
            n_Body_x[739] = c_Body_x[739];
            n_Body_y[739] = c_Body_y[739];
            n_Body_x[740] = c_Body_x[740];
            n_Body_y[740] = c_Body_y[740];
            n_Body_x[741] = c_Body_x[741];
            n_Body_y[741] = c_Body_y[741];
            n_Body_x[742] = c_Body_x[742];
            n_Body_y[742] = c_Body_y[742];
            n_Body_x[743] = c_Body_x[743];
            n_Body_y[743] = c_Body_y[743];
            n_Body_x[744] = c_Body_x[744];
            n_Body_y[744] = c_Body_y[744];
            n_Body_x[745] = c_Body_x[745];
            n_Body_y[745] = c_Body_y[745];
            n_Body_x[746] = c_Body_x[746];
            n_Body_y[746] = c_Body_y[746];
            n_Body_x[747] = c_Body_x[747];
            n_Body_y[747] = c_Body_y[747];
            n_Body_x[748] = c_Body_x[748];
            n_Body_y[748] = c_Body_y[748];
            n_Body_x[749] = c_Body_x[749];
            n_Body_y[749] = c_Body_y[749];
            n_Body_x[750] = c_Body_x[750];
            n_Body_y[750] = c_Body_y[750];
            n_Body_x[751] = c_Body_x[751];
            n_Body_y[751] = c_Body_y[751];
            n_Body_x[752] = c_Body_x[752];
            n_Body_y[752] = c_Body_y[752];
            n_Body_x[753] = c_Body_x[753];
            n_Body_y[753] = c_Body_y[753];
            n_Body_x[754] = c_Body_x[754];
            n_Body_y[754] = c_Body_y[754];
            n_Body_x[755] = c_Body_x[755];
            n_Body_y[755] = c_Body_y[755];
            n_Body_x[756] = c_Body_x[756];
            n_Body_y[756] = c_Body_y[756];
            n_Body_x[757] = c_Body_x[757];
            n_Body_y[757] = c_Body_y[757];
            n_Body_x[758] = c_Body_x[758];
            n_Body_y[758] = c_Body_y[758];
            n_Body_x[759] = c_Body_x[759];
            n_Body_y[759] = c_Body_y[759];
            n_Body_x[760] = c_Body_x[760];
            n_Body_y[760] = c_Body_y[760];
            n_Body_x[761] = c_Body_x[761];
            n_Body_y[761] = c_Body_y[761];
            n_Body_x[762] = c_Body_x[762];
            n_Body_y[762] = c_Body_y[762];
            n_Body_x[763] = c_Body_x[763];
            n_Body_y[763] = c_Body_y[763];
            n_Body_x[764] = c_Body_x[764];
            n_Body_y[764] = c_Body_y[764];
            n_Body_x[765] = c_Body_x[765];
            n_Body_y[765] = c_Body_y[765];
            n_Body_x[766] = c_Body_x[766];
            n_Body_y[766] = c_Body_y[766];
            n_Body_x[767] = c_Body_x[767];
            n_Body_y[767] = c_Body_y[767];
            n_Body_x[768] = c_Body_x[768];
            n_Body_y[768] = c_Body_y[768];
            n_Body_x[769] = c_Body_x[769];
            n_Body_y[769] = c_Body_y[769];
            n_Body_x[770] = c_Body_x[770];
            n_Body_y[770] = c_Body_y[770];
            n_Body_x[771] = c_Body_x[771];
            n_Body_y[771] = c_Body_y[771];
            n_Body_x[772] = c_Body_x[772];
            n_Body_y[772] = c_Body_y[772];
            n_Body_x[773] = c_Body_x[773];
            n_Body_y[773] = c_Body_y[773];
            n_Body_x[774] = c_Body_x[774];
            n_Body_y[774] = c_Body_y[774];
            n_Body_x[775] = c_Body_x[775];
            n_Body_y[775] = c_Body_y[775];
            n_Body_x[776] = c_Body_x[776];
            n_Body_y[776] = c_Body_y[776];
            n_Body_x[777] = c_Body_x[777];
            n_Body_y[777] = c_Body_y[777];
            n_Body_x[778] = c_Body_x[778];
            n_Body_y[778] = c_Body_y[778];
            n_Body_x[779] = c_Body_x[779];
            n_Body_y[779] = c_Body_y[779];
            n_Body_x[780] = c_Body_x[780];
            n_Body_y[780] = c_Body_y[780];
            n_Body_x[781] = c_Body_x[781];
            n_Body_y[781] = c_Body_y[781];
            n_Body_x[782] = c_Body_x[782];
            n_Body_y[782] = c_Body_y[782];
            n_Body_x[783] = c_Body_x[783];
            n_Body_y[783] = c_Body_y[783];
            n_Body_x[784] = c_Body_x[784];
            n_Body_y[784] = c_Body_y[784];
            n_Body_x[785] = c_Body_x[785];
            n_Body_y[785] = c_Body_y[785];
            n_Body_x[786] = c_Body_x[786];
            n_Body_y[786] = c_Body_y[786];
            n_Body_x[787] = c_Body_x[787];
            n_Body_y[787] = c_Body_y[787];
            n_Body_x[788] = c_Body_x[788];
            n_Body_y[788] = c_Body_y[788];
            n_Body_x[789] = c_Body_x[789];
            n_Body_y[789] = c_Body_y[789];
            n_Body_x[790] = c_Body_x[790];
            n_Body_y[790] = c_Body_y[790];
            n_Body_x[791] = c_Body_x[791];
            n_Body_y[791] = c_Body_y[791];
            n_Body_x[792] = c_Body_x[792];
            n_Body_y[792] = c_Body_y[792];
            n_Body_x[793] = c_Body_x[793];
            n_Body_y[793] = c_Body_y[793];
            n_Body_x[794] = c_Body_x[794];
            n_Body_y[794] = c_Body_y[794];
            n_Body_x[795] = c_Body_x[795];
            n_Body_y[795] = c_Body_y[795];
            n_Body_x[796] = c_Body_x[796];
            n_Body_y[796] = c_Body_y[796];
            n_Body_x[797] = c_Body_x[797];
            n_Body_y[797] = c_Body_y[797];
            n_Body_x[798] = c_Body_x[798];
            n_Body_y[798] = c_Body_y[798];
            n_Body_x[799] = c_Body_x[799];
            n_Body_y[799] = c_Body_y[799];
            n_Body_x[800] = c_Body_x[800];
            n_Body_y[800] = c_Body_y[800];
            n_Body_x[801] = c_Body_x[801];
            n_Body_y[801] = c_Body_y[801];
            n_Body_x[802] = c_Body_x[802];
            n_Body_y[802] = c_Body_y[802];
            n_Body_x[803] = c_Body_x[803];
            n_Body_y[803] = c_Body_y[803];
            n_Body_x[804] = c_Body_x[804];
            n_Body_y[804] = c_Body_y[804];
            n_Body_x[805] = c_Body_x[805];
            n_Body_y[805] = c_Body_y[805];
            n_Body_x[806] = c_Body_x[806];
            n_Body_y[806] = c_Body_y[806];
            n_Body_x[807] = c_Body_x[807];
            n_Body_y[807] = c_Body_y[807];
            n_Body_x[808] = c_Body_x[808];
            n_Body_y[808] = c_Body_y[808];
            n_Body_x[809] = c_Body_x[809];
            n_Body_y[809] = c_Body_y[809];
            n_Body_x[810] = c_Body_x[810];
            n_Body_y[810] = c_Body_y[810];
            n_Body_x[811] = c_Body_x[811];
            n_Body_y[811] = c_Body_y[811];
            n_Body_x[812] = c_Body_x[812];
            n_Body_y[812] = c_Body_y[812];
            n_Body_x[813] = c_Body_x[813];
            n_Body_y[813] = c_Body_y[813];
            n_Body_x[814] = c_Body_x[814];
            n_Body_y[814] = c_Body_y[814];
            n_Body_x[815] = c_Body_x[815];
            n_Body_y[815] = c_Body_y[815];
            n_Body_x[816] = c_Body_x[816];
            n_Body_y[816] = c_Body_y[816];
            n_Body_x[817] = c_Body_x[817];
            n_Body_y[817] = c_Body_y[817];
            n_Body_x[818] = c_Body_x[818];
            n_Body_y[818] = c_Body_y[818];
            n_Body_x[819] = c_Body_x[819];
            n_Body_y[819] = c_Body_y[819];
            n_Body_x[820] = c_Body_x[820];
            n_Body_y[820] = c_Body_y[820];
            n_Body_x[821] = c_Body_x[821];
            n_Body_y[821] = c_Body_y[821];
            n_Body_x[822] = c_Body_x[822];
            n_Body_y[822] = c_Body_y[822];
            n_Body_x[823] = c_Body_x[823];
            n_Body_y[823] = c_Body_y[823];
            n_Body_x[824] = c_Body_x[824];
            n_Body_y[824] = c_Body_y[824];
            n_Body_x[825] = c_Body_x[825];
            n_Body_y[825] = c_Body_y[825];
            n_Body_x[826] = c_Body_x[826];
            n_Body_y[826] = c_Body_y[826];
            n_Body_x[827] = c_Body_x[827];
            n_Body_y[827] = c_Body_y[827];
            n_Body_x[828] = c_Body_x[828];
            n_Body_y[828] = c_Body_y[828];
            n_Body_x[829] = c_Body_x[829];
            n_Body_y[829] = c_Body_y[829];
            n_Body_x[830] = c_Body_x[830];
            n_Body_y[830] = c_Body_y[830];
            n_Body_x[831] = c_Body_x[831];
            n_Body_y[831] = c_Body_y[831];
            n_Body_x[832] = c_Body_x[832];
            n_Body_y[832] = c_Body_y[832];
            n_Body_x[833] = c_Body_x[833];
            n_Body_y[833] = c_Body_y[833];
            n_Body_x[834] = c_Body_x[834];
            n_Body_y[834] = c_Body_y[834];
            n_Body_x[835] = c_Body_x[835];
            n_Body_y[835] = c_Body_y[835];
            n_Body_x[836] = c_Body_x[836];
            n_Body_y[836] = c_Body_y[836];
            n_Body_x[837] = c_Body_x[837];
            n_Body_y[837] = c_Body_y[837];
            n_Body_x[838] = c_Body_x[838];
            n_Body_y[838] = c_Body_y[838];
            n_Body_x[839] = c_Body_x[839];
            n_Body_y[839] = c_Body_y[839];
            n_Body_x[840] = c_Body_x[840];
            n_Body_y[840] = c_Body_y[840];
            n_Body_x[841] = c_Body_x[841];
            n_Body_y[841] = c_Body_y[841];
            n_Body_x[842] = c_Body_x[842];
            n_Body_y[842] = c_Body_y[842];
            n_Body_x[843] = c_Body_x[843];
            n_Body_y[843] = c_Body_y[843];
            n_Body_x[844] = c_Body_x[844];
            n_Body_y[844] = c_Body_y[844];
            n_Body_x[845] = c_Body_x[845];
            n_Body_y[845] = c_Body_y[845];
            n_Body_x[846] = c_Body_x[846];
            n_Body_y[846] = c_Body_y[846];
            n_Body_x[847] = c_Body_x[847];
            n_Body_y[847] = c_Body_y[847];
            n_Body_x[848] = c_Body_x[848];
            n_Body_y[848] = c_Body_y[848];
            n_Body_x[849] = c_Body_x[849];
            n_Body_y[849] = c_Body_y[849];
            n_Body_x[850] = c_Body_x[850];
            n_Body_y[850] = c_Body_y[850];
            n_Body_x[851] = c_Body_x[851];
            n_Body_y[851] = c_Body_y[851];
            n_Body_x[852] = c_Body_x[852];
            n_Body_y[852] = c_Body_y[852];
            n_Body_x[853] = c_Body_x[853];
            n_Body_y[853] = c_Body_y[853];
            n_Body_x[854] = c_Body_x[854];
            n_Body_y[854] = c_Body_y[854];
            n_Body_x[855] = c_Body_x[855];
            n_Body_y[855] = c_Body_y[855];
            n_Body_x[856] = c_Body_x[856];
            n_Body_y[856] = c_Body_y[856];
            n_Body_x[857] = c_Body_x[857];
            n_Body_y[857] = c_Body_y[857];
            n_Body_x[858] = c_Body_x[858];
            n_Body_y[858] = c_Body_y[858];
            n_Body_x[859] = c_Body_x[859];
            n_Body_y[859] = c_Body_y[859];
            n_Body_x[860] = c_Body_x[860];
            n_Body_y[860] = c_Body_y[860];
            n_Body_x[861] = c_Body_x[861];
            n_Body_y[861] = c_Body_y[861];
            n_Body_x[862] = c_Body_x[862];
            n_Body_y[862] = c_Body_y[862];
            n_Body_x[863] = c_Body_x[863];
            n_Body_y[863] = c_Body_y[863];
            n_Body_x[864] = c_Body_x[864];
            n_Body_y[864] = c_Body_y[864];
            n_Body_x[865] = c_Body_x[865];
            n_Body_y[865] = c_Body_y[865];
            n_Body_x[866] = c_Body_x[866];
            n_Body_y[866] = c_Body_y[866];
            n_Body_x[867] = c_Body_x[867];
            n_Body_y[867] = c_Body_y[867];
            n_Body_x[868] = c_Body_x[868];
            n_Body_y[868] = c_Body_y[868];
            n_Body_x[869] = c_Body_x[869];
            n_Body_y[869] = c_Body_y[869];
            n_Body_x[870] = c_Body_x[870];
            n_Body_y[870] = c_Body_y[870];
            n_Body_x[871] = c_Body_x[871];
            n_Body_y[871] = c_Body_y[871];
            n_Body_x[872] = c_Body_x[872];
            n_Body_y[872] = c_Body_y[872];
            n_Body_x[873] = c_Body_x[873];
            n_Body_y[873] = c_Body_y[873];
            n_Body_x[874] = c_Body_x[874];
            n_Body_y[874] = c_Body_y[874];
            n_Body_x[875] = c_Body_x[875];
            n_Body_y[875] = c_Body_y[875];
            n_Body_x[876] = c_Body_x[876];
            n_Body_y[876] = c_Body_y[876];
            n_Body_x[877] = c_Body_x[877];
            n_Body_y[877] = c_Body_y[877];
            n_Body_x[878] = c_Body_x[878];
            n_Body_y[878] = c_Body_y[878];
            n_Body_x[879] = c_Body_x[879];
            n_Body_y[879] = c_Body_y[879];
            n_Body_x[880] = c_Body_x[880];
            n_Body_y[880] = c_Body_y[880];
            n_Body_x[881] = c_Body_x[881];
            n_Body_y[881] = c_Body_y[881];
            n_Body_x[882] = c_Body_x[882];
            n_Body_y[882] = c_Body_y[882];
            n_Body_x[883] = c_Body_x[883];
            n_Body_y[883] = c_Body_y[883];
            n_Body_x[884] = c_Body_x[884];
            n_Body_y[884] = c_Body_y[884];
            n_Body_x[885] = c_Body_x[885];
            n_Body_y[885] = c_Body_y[885];
            n_Body_x[886] = c_Body_x[886];
            n_Body_y[886] = c_Body_y[886];
            n_Body_x[887] = c_Body_x[887];
            n_Body_y[887] = c_Body_y[887];
            n_Body_x[888] = c_Body_x[888];
            n_Body_y[888] = c_Body_y[888];
            n_Body_x[889] = c_Body_x[889];
            n_Body_y[889] = c_Body_y[889];
            n_Body_x[890] = c_Body_x[890];
            n_Body_y[890] = c_Body_y[890];
            n_Body_x[891] = c_Body_x[891];
            n_Body_y[891] = c_Body_y[891];
            n_Body_x[892] = c_Body_x[892];
            n_Body_y[892] = c_Body_y[892];
            n_Body_x[893] = c_Body_x[893];
            n_Body_y[893] = c_Body_y[893];
            n_Body_x[894] = c_Body_x[894];
            n_Body_y[894] = c_Body_y[894];
            n_Body_x[895] = c_Body_x[895];
            n_Body_y[895] = c_Body_y[895];
            n_Body_x[896] = c_Body_x[896];
            n_Body_y[896] = c_Body_y[896];
            n_Body_x[897] = c_Body_x[897];
            n_Body_y[897] = c_Body_y[897];
            n_Body_x[898] = c_Body_x[898];
            n_Body_y[898] = c_Body_y[898];
            n_Body_x[899] = c_Body_x[899];
            n_Body_y[899] = c_Body_y[899];
            n_Body_x[900] = c_Body_x[900];
            n_Body_y[900] = c_Body_y[900];
            n_Body_x[901] = c_Body_x[901];
            n_Body_y[901] = c_Body_y[901];
            n_Body_x[902] = c_Body_x[902];
            n_Body_y[902] = c_Body_y[902];
            n_Body_x[903] = c_Body_x[903];
            n_Body_y[903] = c_Body_y[903];
            n_Body_x[904] = c_Body_x[904];
            n_Body_y[904] = c_Body_y[904];
            n_Body_x[905] = c_Body_x[905];
            n_Body_y[905] = c_Body_y[905];
            n_Body_x[906] = c_Body_x[906];
            n_Body_y[906] = c_Body_y[906];
            n_Body_x[907] = c_Body_x[907];
            n_Body_y[907] = c_Body_y[907];
            n_Body_x[908] = c_Body_x[908];
            n_Body_y[908] = c_Body_y[908];
            n_Body_x[909] = c_Body_x[909];
            n_Body_y[909] = c_Body_y[909];
            n_Body_x[910] = c_Body_x[910];
            n_Body_y[910] = c_Body_y[910];
            n_Body_x[911] = c_Body_x[911];
            n_Body_y[911] = c_Body_y[911];
            n_Body_x[912] = c_Body_x[912];
            n_Body_y[912] = c_Body_y[912];
            n_Body_x[913] = c_Body_x[913];
            n_Body_y[913] = c_Body_y[913];
            n_Body_x[914] = c_Body_x[914];
            n_Body_y[914] = c_Body_y[914];
            n_Body_x[915] = c_Body_x[915];
            n_Body_y[915] = c_Body_y[915];
            n_Body_x[916] = c_Body_x[916];
            n_Body_y[916] = c_Body_y[916];
            n_Body_x[917] = c_Body_x[917];
            n_Body_y[917] = c_Body_y[917];
            n_Body_x[918] = c_Body_x[918];
            n_Body_y[918] = c_Body_y[918];
            n_Body_x[919] = c_Body_x[919];
            n_Body_y[919] = c_Body_y[919];
            n_Body_x[920] = c_Body_x[920];
            n_Body_y[920] = c_Body_y[920];
            n_Body_x[921] = c_Body_x[921];
            n_Body_y[921] = c_Body_y[921];
            n_Body_x[922] = c_Body_x[922];
            n_Body_y[922] = c_Body_y[922];
            n_Body_x[923] = c_Body_x[923];
            n_Body_y[923] = c_Body_y[923];
            n_Body_x[924] = c_Body_x[924];
            n_Body_y[924] = c_Body_y[924];
            n_Body_x[925] = c_Body_x[925];
            n_Body_y[925] = c_Body_y[925];
            n_Body_x[926] = c_Body_x[926];
            n_Body_y[926] = c_Body_y[926];
            n_Body_x[927] = c_Body_x[927];
            n_Body_y[927] = c_Body_y[927];
            n_Body_x[928] = c_Body_x[928];
            n_Body_y[928] = c_Body_y[928];
            n_Body_x[929] = c_Body_x[929];
            n_Body_y[929] = c_Body_y[929];
            n_Body_x[930] = c_Body_x[930];
            n_Body_y[930] = c_Body_y[930];
            n_Body_x[931] = c_Body_x[931];
            n_Body_y[931] = c_Body_y[931];
            n_Body_x[932] = c_Body_x[932];
            n_Body_y[932] = c_Body_y[932];
            n_Body_x[933] = c_Body_x[933];
            n_Body_y[933] = c_Body_y[933];
            n_Body_x[934] = c_Body_x[934];
            n_Body_y[934] = c_Body_y[934];
            n_Body_x[935] = c_Body_x[935];
            n_Body_y[935] = c_Body_y[935];
            n_Body_x[936] = c_Body_x[936];
            n_Body_y[936] = c_Body_y[936];
            n_Body_x[937] = c_Body_x[937];
            n_Body_y[937] = c_Body_y[937];
            n_Body_x[938] = c_Body_x[938];
            n_Body_y[938] = c_Body_y[938];
            n_Body_x[939] = c_Body_x[939];
            n_Body_y[939] = c_Body_y[939];
            n_Body_x[940] = c_Body_x[940];
            n_Body_y[940] = c_Body_y[940];
            n_Body_x[941] = c_Body_x[941];
            n_Body_y[941] = c_Body_y[941];
            n_Body_x[942] = c_Body_x[942];
            n_Body_y[942] = c_Body_y[942];
            n_Body_x[943] = c_Body_x[943];
            n_Body_y[943] = c_Body_y[943];
            n_Body_x[944] = c_Body_x[944];
            n_Body_y[944] = c_Body_y[944];
            n_Body_x[945] = c_Body_x[945];
            n_Body_y[945] = c_Body_y[945];
            n_Body_x[946] = c_Body_x[946];
            n_Body_y[946] = c_Body_y[946];
            n_Body_x[947] = c_Body_x[947];
            n_Body_y[947] = c_Body_y[947];
            n_Body_x[948] = c_Body_x[948];
            n_Body_y[948] = c_Body_y[948];
            n_Body_x[949] = c_Body_x[949];
            n_Body_y[949] = c_Body_y[949];
            n_Body_x[950] = c_Body_x[950];
            n_Body_y[950] = c_Body_y[950];
            n_Body_x[951] = c_Body_x[951];
            n_Body_y[951] = c_Body_y[951];
            n_Body_x[952] = c_Body_x[952];
            n_Body_y[952] = c_Body_y[952];
            n_Body_x[953] = c_Body_x[953];
            n_Body_y[953] = c_Body_y[953];
            n_Body_x[954] = c_Body_x[954];
            n_Body_y[954] = c_Body_y[954];
            n_Body_x[955] = c_Body_x[955];
            n_Body_y[955] = c_Body_y[955];
            n_Body_x[956] = c_Body_x[956];
            n_Body_y[956] = c_Body_y[956];
            n_Body_x[957] = c_Body_x[957];
            n_Body_y[957] = c_Body_y[957];
            n_Body_x[958] = c_Body_x[958];
            n_Body_y[958] = c_Body_y[958];
            n_Body_x[959] = c_Body_x[959];
            n_Body_y[959] = c_Body_y[959];
            n_Body_x[960] = c_Body_x[960];
            n_Body_y[960] = c_Body_y[960];
            n_Body_x[961] = c_Body_x[961];
            n_Body_y[961] = c_Body_y[961];
            n_Body_x[962] = c_Body_x[962];
            n_Body_y[962] = c_Body_y[962];
            n_Body_x[963] = c_Body_x[963];
            n_Body_y[963] = c_Body_y[963];
            n_Body_x[964] = c_Body_x[964];
            n_Body_y[964] = c_Body_y[964];
            n_Body_x[965] = c_Body_x[965];
            n_Body_y[965] = c_Body_y[965];
            n_Body_x[966] = c_Body_x[966];
            n_Body_y[966] = c_Body_y[966];
            n_Body_x[967] = c_Body_x[967];
            n_Body_y[967] = c_Body_y[967];
            n_Body_x[968] = c_Body_x[968];
            n_Body_y[968] = c_Body_y[968];
            n_Body_x[969] = c_Body_x[969];
            n_Body_y[969] = c_Body_y[969];
            n_Body_x[970] = c_Body_x[970];
            n_Body_y[970] = c_Body_y[970];
            n_Body_x[971] = c_Body_x[971];
            n_Body_y[971] = c_Body_y[971];
            n_Body_x[972] = c_Body_x[972];
            n_Body_y[972] = c_Body_y[972];
            n_Body_x[973] = c_Body_x[973];
            n_Body_y[973] = c_Body_y[973];
            n_Body_x[974] = c_Body_x[974];
            n_Body_y[974] = c_Body_y[974];
            n_Body_x[975] = c_Body_x[975];
            n_Body_y[975] = c_Body_y[975];
            n_Body_x[976] = c_Body_x[976];
            n_Body_y[976] = c_Body_y[976];
            n_Body_x[977] = c_Body_x[977];
            n_Body_y[977] = c_Body_y[977];
            n_Body_x[978] = c_Body_x[978];
            n_Body_y[978] = c_Body_y[978];
            n_Body_x[979] = c_Body_x[979];
            n_Body_y[979] = c_Body_y[979];
            n_Body_x[980] = c_Body_x[980];
            n_Body_y[980] = c_Body_y[980];
            n_Body_x[981] = c_Body_x[981];
            n_Body_y[981] = c_Body_y[981];
            n_Body_x[982] = c_Body_x[982];
            n_Body_y[982] = c_Body_y[982];
            n_Body_x[983] = c_Body_x[983];
            n_Body_y[983] = c_Body_y[983];
            n_Body_x[984] = c_Body_x[984];
            n_Body_y[984] = c_Body_y[984];
            n_Body_x[985] = c_Body_x[985];
            n_Body_y[985] = c_Body_y[985];
            n_Body_x[986] = c_Body_x[986];
            n_Body_y[986] = c_Body_y[986];
            n_Body_x[987] = c_Body_x[987];
            n_Body_y[987] = c_Body_y[987];
            n_Body_x[988] = c_Body_x[988];
            n_Body_y[988] = c_Body_y[988];
            n_Body_x[989] = c_Body_x[989];
            n_Body_y[989] = c_Body_y[989];
            n_Body_x[990] = c_Body_x[990];
            n_Body_y[990] = c_Body_y[990];
            n_Body_x[991] = c_Body_x[991];
            n_Body_y[991] = c_Body_y[991];
            n_Body_x[992] = c_Body_x[992];
            n_Body_y[992] = c_Body_y[992];
            n_Body_x[993] = c_Body_x[993];
            n_Body_y[993] = c_Body_y[993];
            n_Body_x[994] = c_Body_x[994];
            n_Body_y[994] = c_Body_y[994];
            n_Body_x[995] = c_Body_x[995];
            n_Body_y[995] = c_Body_y[995];
            n_Body_x[996] = c_Body_x[996];
            n_Body_y[996] = c_Body_y[996];
            n_Body_x[997] = c_Body_x[997];
            n_Body_y[997] = c_Body_y[997];
            n_Body_x[998] = c_Body_x[998];
            n_Body_y[998] = c_Body_y[998];
            n_Body_x[999] = c_Body_x[999];
            n_Body_y[999] = c_Body_y[999];
            n_Body_x[1000] = c_Body_x[1000];
            n_Body_y[1000] = c_Body_y[1000];
            n_Body_x[1001] = c_Body_x[1001];
            n_Body_y[1001] = c_Body_y[1001];
            n_Body_x[1002] = c_Body_x[1002];
            n_Body_y[1002] = c_Body_y[1002];
            n_Body_x[1003] = c_Body_x[1003];
            n_Body_y[1003] = c_Body_y[1003];
            n_Body_x[1004] = c_Body_x[1004];
            n_Body_y[1004] = c_Body_y[1004];
            n_Body_x[1005] = c_Body_x[1005];
            n_Body_y[1005] = c_Body_y[1005];
            n_Body_x[1006] = c_Body_x[1006];
            n_Body_y[1006] = c_Body_y[1006];
            n_Body_x[1007] = c_Body_x[1007];
            n_Body_y[1007] = c_Body_y[1007];
            n_Body_x[1008] = c_Body_x[1008];
            n_Body_y[1008] = c_Body_y[1008];
            n_Body_x[1009] = c_Body_x[1009];
            n_Body_y[1009] = c_Body_y[1009];
            n_Body_x[1010] = c_Body_x[1010];
            n_Body_y[1010] = c_Body_y[1010];
            n_Body_x[1011] = c_Body_x[1011];
            n_Body_y[1011] = c_Body_y[1011];
            n_Body_x[1012] = c_Body_x[1012];
            n_Body_y[1012] = c_Body_y[1012];
            n_Body_x[1013] = c_Body_x[1013];
            n_Body_y[1013] = c_Body_y[1013];
            n_Body_x[1014] = c_Body_x[1014];
            n_Body_y[1014] = c_Body_y[1014];
            n_Body_x[1015] = c_Body_x[1015];
            n_Body_y[1015] = c_Body_y[1015];
            n_Body_x[1016] = c_Body_x[1016];
            n_Body_y[1016] = c_Body_y[1016];
            n_Body_x[1017] = c_Body_x[1017];
            n_Body_y[1017] = c_Body_y[1017];
            n_Body_x[1018] = c_Body_x[1018];
            n_Body_y[1018] = c_Body_y[1018];
            n_Body_x[1019] = c_Body_x[1019];
            n_Body_y[1019] = c_Body_y[1019];
            n_Body_x[1020] = c_Body_x[1020];
            n_Body_y[1020] = c_Body_y[1020];
            n_Body_x[1021] = c_Body_x[1021];
            n_Body_y[1021] = c_Body_y[1021];
            n_Body_x[1022] = c_Body_x[1022];
            n_Body_y[1022] = c_Body_y[1022];
            n_Body_x[1023] = c_Body_x[1023];
            n_Body_y[1023] = c_Body_y[1023];
            n_Body_x[1024] = c_Body_x[1024];
            n_Body_y[1024] = c_Body_y[1024];
            n_Body_x[1025] = c_Body_x[1025];
            n_Body_y[1025] = c_Body_y[1025];
            n_Body_x[1026] = c_Body_x[1026];
            n_Body_y[1026] = c_Body_y[1026];
            n_Body_x[1027] = c_Body_x[1027];
            n_Body_y[1027] = c_Body_y[1027];
            n_Body_x[1028] = c_Body_x[1028];
            n_Body_y[1028] = c_Body_y[1028];
            n_Body_x[1029] = c_Body_x[1029];
            n_Body_y[1029] = c_Body_y[1029];
            n_Body_x[1030] = c_Body_x[1030];
            n_Body_y[1030] = c_Body_y[1030];
            n_Body_x[1031] = c_Body_x[1031];
            n_Body_y[1031] = c_Body_y[1031];
            n_Body_x[1032] = c_Body_x[1032];
            n_Body_y[1032] = c_Body_y[1032];
            n_Body_x[1033] = c_Body_x[1033];
            n_Body_y[1033] = c_Body_y[1033];
            n_Body_x[1034] = c_Body_x[1034];
            n_Body_y[1034] = c_Body_y[1034];
            n_Body_x[1035] = c_Body_x[1035];
            n_Body_y[1035] = c_Body_y[1035];
            n_Body_x[1036] = c_Body_x[1036];
            n_Body_y[1036] = c_Body_y[1036];
            n_Body_x[1037] = c_Body_x[1037];
            n_Body_y[1037] = c_Body_y[1037];
            n_Body_x[1038] = c_Body_x[1038];
            n_Body_y[1038] = c_Body_y[1038];
            n_Body_x[1039] = c_Body_x[1039];
            n_Body_y[1039] = c_Body_y[1039];
            n_Body_x[1040] = c_Body_x[1040];
            n_Body_y[1040] = c_Body_y[1040];
            n_Body_x[1041] = c_Body_x[1041];
            n_Body_y[1041] = c_Body_y[1041];
            n_Body_x[1042] = c_Body_x[1042];
            n_Body_y[1042] = c_Body_y[1042];
            n_Body_x[1043] = c_Body_x[1043];
            n_Body_y[1043] = c_Body_y[1043];
            n_Body_x[1044] = c_Body_x[1044];
            n_Body_y[1044] = c_Body_y[1044];
            n_Body_x[1045] = c_Body_x[1045];
            n_Body_y[1045] = c_Body_y[1045];
            n_Body_x[1046] = c_Body_x[1046];
            n_Body_y[1046] = c_Body_y[1046];
            n_Body_x[1047] = c_Body_x[1047];
            n_Body_y[1047] = c_Body_y[1047];
            n_Body_x[1048] = c_Body_x[1048];
            n_Body_y[1048] = c_Body_y[1048];
            n_Body_x[1049] = c_Body_x[1049];
            n_Body_y[1049] = c_Body_y[1049];
            n_Body_x[1050] = c_Body_x[1050];
            n_Body_y[1050] = c_Body_y[1050];
            n_Body_x[1051] = c_Body_x[1051];
            n_Body_y[1051] = c_Body_y[1051];
            n_Body_x[1052] = c_Body_x[1052];
            n_Body_y[1052] = c_Body_y[1052];
            n_Body_x[1053] = c_Body_x[1053];
            n_Body_y[1053] = c_Body_y[1053];
            n_Body_x[1054] = c_Body_x[1054];
            n_Body_y[1054] = c_Body_y[1054];
            n_Body_x[1055] = c_Body_x[1055];
            n_Body_y[1055] = c_Body_y[1055];
            n_Body_x[1056] = c_Body_x[1056];
            n_Body_y[1056] = c_Body_y[1056];
            n_Body_x[1057] = c_Body_x[1057];
            n_Body_y[1057] = c_Body_y[1057];
            n_Body_x[1058] = c_Body_x[1058];
            n_Body_y[1058] = c_Body_y[1058];
            n_Body_x[1059] = c_Body_x[1059];
            n_Body_y[1059] = c_Body_y[1059];
            n_Body_x[1060] = c_Body_x[1060];
            n_Body_y[1060] = c_Body_y[1060];
            n_Body_x[1061] = c_Body_x[1061];
            n_Body_y[1061] = c_Body_y[1061];
            n_Body_x[1062] = c_Body_x[1062];
            n_Body_y[1062] = c_Body_y[1062];
            n_Body_x[1063] = c_Body_x[1063];
            n_Body_y[1063] = c_Body_y[1063];
            n_Body_x[1064] = c_Body_x[1064];
            n_Body_y[1064] = c_Body_y[1064];
            n_Body_x[1065] = c_Body_x[1065];
            n_Body_y[1065] = c_Body_y[1065];
            n_Body_x[1066] = c_Body_x[1066];
            n_Body_y[1066] = c_Body_y[1066];
            n_Body_x[1067] = c_Body_x[1067];
            n_Body_y[1067] = c_Body_y[1067];
            n_Body_x[1068] = c_Body_x[1068];
            n_Body_y[1068] = c_Body_y[1068];
            n_Body_x[1069] = c_Body_x[1069];
            n_Body_y[1069] = c_Body_y[1069];
            n_Body_x[1070] = c_Body_x[1070];
            n_Body_y[1070] = c_Body_y[1070];
            n_Body_x[1071] = c_Body_x[1071];
            n_Body_y[1071] = c_Body_y[1071];
            n_Body_x[1072] = c_Body_x[1072];
            n_Body_y[1072] = c_Body_y[1072];
            n_Body_x[1073] = c_Body_x[1073];
            n_Body_y[1073] = c_Body_y[1073];
            n_Body_x[1074] = c_Body_x[1074];
            n_Body_y[1074] = c_Body_y[1074];
            n_Body_x[1075] = c_Body_x[1075];
            n_Body_y[1075] = c_Body_y[1075];
            n_Body_x[1076] = c_Body_x[1076];
            n_Body_y[1076] = c_Body_y[1076];
            n_Body_x[1077] = c_Body_x[1077];
            n_Body_y[1077] = c_Body_y[1077];
            n_Body_x[1078] = c_Body_x[1078];
            n_Body_y[1078] = c_Body_y[1078];
            n_Body_x[1079] = c_Body_x[1079];
            n_Body_y[1079] = c_Body_y[1079];
            n_Body_x[1080] = c_Body_x[1080];
            n_Body_y[1080] = c_Body_y[1080];
            n_Body_x[1081] = c_Body_x[1081];
            n_Body_y[1081] = c_Body_y[1081];
            n_Body_x[1082] = c_Body_x[1082];
            n_Body_y[1082] = c_Body_y[1082];
            n_Body_x[1083] = c_Body_x[1083];
            n_Body_y[1083] = c_Body_y[1083];
            n_Body_x[1084] = c_Body_x[1084];
            n_Body_y[1084] = c_Body_y[1084];
            n_Body_x[1085] = c_Body_x[1085];
            n_Body_y[1085] = c_Body_y[1085];
            n_Body_x[1086] = c_Body_x[1086];
            n_Body_y[1086] = c_Body_y[1086];
            n_Body_x[1087] = c_Body_x[1087];
            n_Body_y[1087] = c_Body_y[1087];
            n_Body_x[1088] = c_Body_x[1088];
            n_Body_y[1088] = c_Body_y[1088];
            n_Body_x[1089] = c_Body_x[1089];
            n_Body_y[1089] = c_Body_y[1089];
            n_Body_x[1090] = c_Body_x[1090];
            n_Body_y[1090] = c_Body_y[1090];
            n_Body_x[1091] = c_Body_x[1091];
            n_Body_y[1091] = c_Body_y[1091];
            n_Body_x[1092] = c_Body_x[1092];
            n_Body_y[1092] = c_Body_y[1092];
            n_Body_x[1093] = c_Body_x[1093];
            n_Body_y[1093] = c_Body_y[1093];
            n_Body_x[1094] = c_Body_x[1094];
            n_Body_y[1094] = c_Body_y[1094];
            n_Body_x[1095] = c_Body_x[1095];
            n_Body_y[1095] = c_Body_y[1095];
            n_Body_x[1096] = c_Body_x[1096];
            n_Body_y[1096] = c_Body_y[1096];
            n_Body_x[1097] = c_Body_x[1097];
            n_Body_y[1097] = c_Body_y[1097];
            n_Body_x[1098] = c_Body_x[1098];
            n_Body_y[1098] = c_Body_y[1098];
            n_Body_x[1099] = c_Body_x[1099];
            n_Body_y[1099] = c_Body_y[1099];
            n_Body_x[1100] = c_Body_x[1100];
            n_Body_y[1100] = c_Body_y[1100];
            n_Body_x[1101] = c_Body_x[1101];
            n_Body_y[1101] = c_Body_y[1101];
            n_Body_x[1102] = c_Body_x[1102];
            n_Body_y[1102] = c_Body_y[1102];
            n_Body_x[1103] = c_Body_x[1103];
            n_Body_y[1103] = c_Body_y[1103];
            n_Body_x[1104] = c_Body_x[1104];
            n_Body_y[1104] = c_Body_y[1104];
            n_Body_x[1105] = c_Body_x[1105];
            n_Body_y[1105] = c_Body_y[1105];
            n_Body_x[1106] = c_Body_x[1106];
            n_Body_y[1106] = c_Body_y[1106];
            n_Body_x[1107] = c_Body_x[1107];
            n_Body_y[1107] = c_Body_y[1107];
            n_Body_x[1108] = c_Body_x[1108];
            n_Body_y[1108] = c_Body_y[1108];
            n_Body_x[1109] = c_Body_x[1109];
            n_Body_y[1109] = c_Body_y[1109];
            n_Body_x[1110] = c_Body_x[1110];
            n_Body_y[1110] = c_Body_y[1110];
            n_Body_x[1111] = c_Body_x[1111];
            n_Body_y[1111] = c_Body_y[1111];
            n_Body_x[1112] = c_Body_x[1112];
            n_Body_y[1112] = c_Body_y[1112];
            n_Body_x[1113] = c_Body_x[1113];
            n_Body_y[1113] = c_Body_y[1113];
            n_Body_x[1114] = c_Body_x[1114];
            n_Body_y[1114] = c_Body_y[1114];
            n_Body_x[1115] = c_Body_x[1115];
            n_Body_y[1115] = c_Body_y[1115];
            n_Body_x[1116] = c_Body_x[1116];
            n_Body_y[1116] = c_Body_y[1116];
            n_Body_x[1117] = c_Body_x[1117];
            n_Body_y[1117] = c_Body_y[1117];
            n_Body_x[1118] = c_Body_x[1118];
            n_Body_y[1118] = c_Body_y[1118];
            n_Body_x[1119] = c_Body_x[1119];
            n_Body_y[1119] = c_Body_y[1119];
            n_Body_x[1120] = c_Body_x[1120];
            n_Body_y[1120] = c_Body_y[1120];
            n_Body_x[1121] = c_Body_x[1121];
            n_Body_y[1121] = c_Body_y[1121];
            n_Body_x[1122] = c_Body_x[1122];
            n_Body_y[1122] = c_Body_y[1122];
            n_Body_x[1123] = c_Body_x[1123];
            n_Body_y[1123] = c_Body_y[1123];
            n_Body_x[1124] = c_Body_x[1124];
            n_Body_y[1124] = c_Body_y[1124];
            n_Body_x[1125] = c_Body_x[1125];
            n_Body_y[1125] = c_Body_y[1125];
            n_Body_x[1126] = c_Body_x[1126];
            n_Body_y[1126] = c_Body_y[1126];
            n_Body_x[1127] = c_Body_x[1127];
            n_Body_y[1127] = c_Body_y[1127];
            n_Body_x[1128] = c_Body_x[1128];
            n_Body_y[1128] = c_Body_y[1128];
            n_Body_x[1129] = c_Body_x[1129];
            n_Body_y[1129] = c_Body_y[1129];
            n_Body_x[1130] = c_Body_x[1130];
            n_Body_y[1130] = c_Body_y[1130];
            n_Body_x[1131] = c_Body_x[1131];
            n_Body_y[1131] = c_Body_y[1131];
            n_Body_x[1132] = c_Body_x[1132];
            n_Body_y[1132] = c_Body_y[1132];
            n_Body_x[1133] = c_Body_x[1133];
            n_Body_y[1133] = c_Body_y[1133];
            n_Body_x[1134] = c_Body_x[1134];
            n_Body_y[1134] = c_Body_y[1134];
            n_Body_x[1135] = c_Body_x[1135];
            n_Body_y[1135] = c_Body_y[1135];
            n_Body_x[1136] = c_Body_x[1136];
            n_Body_y[1136] = c_Body_y[1136];
            n_Body_x[1137] = c_Body_x[1137];
            n_Body_y[1137] = c_Body_y[1137];
            n_Body_x[1138] = c_Body_x[1138];
            n_Body_y[1138] = c_Body_y[1138];
            n_Body_x[1139] = c_Body_x[1139];
            n_Body_y[1139] = c_Body_y[1139];
            n_Body_x[1140] = c_Body_x[1140];
            n_Body_y[1140] = c_Body_y[1140];
            n_Body_x[1141] = c_Body_x[1141];
            n_Body_y[1141] = c_Body_y[1141];
            n_Body_x[1142] = c_Body_x[1142];
            n_Body_y[1142] = c_Body_y[1142];
            n_Body_x[1143] = c_Body_x[1143];
            n_Body_y[1143] = c_Body_y[1143];
            n_Body_x[1144] = c_Body_x[1144];
            n_Body_y[1144] = c_Body_y[1144];
            n_Body_x[1145] = c_Body_x[1145];
            n_Body_y[1145] = c_Body_y[1145];
            n_Body_x[1146] = c_Body_x[1146];
            n_Body_y[1146] = c_Body_y[1146];
            n_Body_x[1147] = c_Body_x[1147];
            n_Body_y[1147] = c_Body_y[1147];
            n_Body_x[1148] = c_Body_x[1148];
            n_Body_y[1148] = c_Body_y[1148];
            n_Body_x[1149] = c_Body_x[1149];
            n_Body_y[1149] = c_Body_y[1149];
            n_Body_x[1150] = c_Body_x[1150];
            n_Body_y[1150] = c_Body_y[1150];
            n_Body_x[1151] = c_Body_x[1151];
            n_Body_y[1151] = c_Body_y[1151];
            n_Body_x[1152] = c_Body_x[1152];
            n_Body_y[1152] = c_Body_y[1152];
            n_Body_x[1153] = c_Body_x[1153];
            n_Body_y[1153] = c_Body_y[1153];
            n_Body_x[1154] = c_Body_x[1154];
            n_Body_y[1154] = c_Body_y[1154];
            n_Body_x[1155] = c_Body_x[1155];
            n_Body_y[1155] = c_Body_y[1155];
            n_Body_x[1156] = c_Body_x[1156];
            n_Body_y[1156] = c_Body_y[1156];
            n_Body_x[1157] = c_Body_x[1157];
            n_Body_y[1157] = c_Body_y[1157];
            n_Body_x[1158] = c_Body_x[1158];
            n_Body_y[1158] = c_Body_y[1158];
            n_Body_x[1159] = c_Body_x[1159];
            n_Body_y[1159] = c_Body_y[1159];
            n_Body_x[1160] = c_Body_x[1160];
            n_Body_y[1160] = c_Body_y[1160];
            n_Body_x[1161] = c_Body_x[1161];
            n_Body_y[1161] = c_Body_y[1161];
            n_Body_x[1162] = c_Body_x[1162];
            n_Body_y[1162] = c_Body_y[1162];
            n_Body_x[1163] = c_Body_x[1163];
            n_Body_y[1163] = c_Body_y[1163];
            n_Body_x[1164] = c_Body_x[1164];
            n_Body_y[1164] = c_Body_y[1164];
            n_Body_x[1165] = c_Body_x[1165];
            n_Body_y[1165] = c_Body_y[1165];
            n_Body_x[1166] = c_Body_x[1166];
            n_Body_y[1166] = c_Body_y[1166];
            n_Body_x[1167] = c_Body_x[1167];
            n_Body_y[1167] = c_Body_y[1167];
            n_Body_x[1168] = c_Body_x[1168];
            n_Body_y[1168] = c_Body_y[1168];
            n_Body_x[1169] = c_Body_x[1169];
            n_Body_y[1169] = c_Body_y[1169];
            n_Body_x[1170] = c_Body_x[1170];
            n_Body_y[1170] = c_Body_y[1170];
            n_Body_x[1171] = c_Body_x[1171];
            n_Body_y[1171] = c_Body_y[1171];
            n_Body_x[1172] = c_Body_x[1172];
            n_Body_y[1172] = c_Body_y[1172];
            n_Body_x[1173] = c_Body_x[1173];
            n_Body_y[1173] = c_Body_y[1173];
            n_Body_x[1174] = c_Body_x[1174];
            n_Body_y[1174] = c_Body_y[1174];
            n_Body_x[1175] = c_Body_x[1175];
            n_Body_y[1175] = c_Body_y[1175];
            n_Body_x[1176] = c_Body_x[1176];
            n_Body_y[1176] = c_Body_y[1176];
            n_Body_x[1177] = c_Body_x[1177];
            n_Body_y[1177] = c_Body_y[1177];
            n_Body_x[1178] = c_Body_x[1178];
            n_Body_y[1178] = c_Body_y[1178];
            n_Body_x[1179] = c_Body_x[1179];
            n_Body_y[1179] = c_Body_y[1179];
            n_Body_x[1180] = c_Body_x[1180];
            n_Body_y[1180] = c_Body_y[1180];
            n_Body_x[1181] = c_Body_x[1181];
            n_Body_y[1181] = c_Body_y[1181];
            n_Body_x[1182] = c_Body_x[1182];
            n_Body_y[1182] = c_Body_y[1182];
            n_Body_x[1183] = c_Body_x[1183];
            n_Body_y[1183] = c_Body_y[1183];
            n_Body_x[1184] = c_Body_x[1184];
            n_Body_y[1184] = c_Body_y[1184];
            n_Body_x[1185] = c_Body_x[1185];
            n_Body_y[1185] = c_Body_y[1185];
            n_Body_x[1186] = c_Body_x[1186];
            n_Body_y[1186] = c_Body_y[1186];
            n_Body_x[1187] = c_Body_x[1187];
            n_Body_y[1187] = c_Body_y[1187];
            n_Body_x[1188] = c_Body_x[1188];
            n_Body_y[1188] = c_Body_y[1188];
            n_Body_x[1189] = c_Body_x[1189];
            n_Body_y[1189] = c_Body_y[1189];
            n_Body_x[1190] = c_Body_x[1190];
            n_Body_y[1190] = c_Body_y[1190];
            n_Body_x[1191] = c_Body_x[1191];
            n_Body_y[1191] = c_Body_y[1191];
            n_Body_x[1192] = c_Body_x[1192];
            n_Body_y[1192] = c_Body_y[1192];
            n_Body_x[1193] = c_Body_x[1193];
            n_Body_y[1193] = c_Body_y[1193];
            n_Body_x[1194] = c_Body_x[1194];
            n_Body_y[1194] = c_Body_y[1194];
            n_Body_x[1195] = c_Body_x[1195];
            n_Body_y[1195] = c_Body_y[1195];
            n_Body_x[1196] = c_Body_x[1196];
            n_Body_y[1196] = c_Body_y[1196];
            n_Body_x[1197] = c_Body_x[1197];
            n_Body_y[1197] = c_Body_y[1197];
            n_Body_x[1198] = c_Body_x[1198];
            n_Body_y[1198] = c_Body_y[1198];
            n_Body_x[1199] = c_Body_x[1199];
            n_Body_y[1199] = c_Body_y[1199];
            n_Body_x[1200] = c_Body_x[1200];
            n_Body_y[1200] = c_Body_y[1200];
            n_Body_x[1201] = c_Body_x[1201];
            n_Body_y[1201] = c_Body_y[1201];
            n_Body_x[1202] = c_Body_x[1202];
            n_Body_y[1202] = c_Body_y[1202];
            n_Body_x[1203] = c_Body_x[1203];
            n_Body_y[1203] = c_Body_y[1203];
            n_Body_x[1204] = c_Body_x[1204];
            n_Body_y[1204] = c_Body_y[1204];
            n_Body_x[1205] = c_Body_x[1205];
            n_Body_y[1205] = c_Body_y[1205];
            n_Body_x[1206] = c_Body_x[1206];
            n_Body_y[1206] = c_Body_y[1206];
            n_Body_x[1207] = c_Body_x[1207];
            n_Body_y[1207] = c_Body_y[1207];
            n_Body_x[1208] = c_Body_x[1208];
            n_Body_y[1208] = c_Body_y[1208];
            n_Body_x[1209] = c_Body_x[1209];
            n_Body_y[1209] = c_Body_y[1209];
            n_Body_x[1210] = c_Body_x[1210];
            n_Body_y[1210] = c_Body_y[1210];
            n_Body_x[1211] = c_Body_x[1211];
            n_Body_y[1211] = c_Body_y[1211];
            n_Body_x[1212] = c_Body_x[1212];
            n_Body_y[1212] = c_Body_y[1212];
            n_Body_x[1213] = c_Body_x[1213];
            n_Body_y[1213] = c_Body_y[1213];
            n_Body_x[1214] = c_Body_x[1214];
            n_Body_y[1214] = c_Body_y[1214];
            n_Body_x[1215] = c_Body_x[1215];
            n_Body_y[1215] = c_Body_y[1215];
            n_Body_x[1216] = c_Body_x[1216];
            n_Body_y[1216] = c_Body_y[1216];
            n_Body_x[1217] = c_Body_x[1217];
            n_Body_y[1217] = c_Body_y[1217];
            n_Body_x[1218] = c_Body_x[1218];
            n_Body_y[1218] = c_Body_y[1218];
            n_Body_x[1219] = c_Body_x[1219];
            n_Body_y[1219] = c_Body_y[1219];
            n_Body_x[1220] = c_Body_x[1220];
            n_Body_y[1220] = c_Body_y[1220];
            n_Body_x[1221] = c_Body_x[1221];
            n_Body_y[1221] = c_Body_y[1221];
            n_Body_x[1222] = c_Body_x[1222];
            n_Body_y[1222] = c_Body_y[1222];
            n_Body_x[1223] = c_Body_x[1223];
            n_Body_y[1223] = c_Body_y[1223];
            n_Body_x[1224] = c_Body_x[1224];
            n_Body_y[1224] = c_Body_y[1224];
            n_Body_x[1225] = c_Body_x[1225];
            n_Body_y[1225] = c_Body_y[1225];
            n_Body_x[1226] = c_Body_x[1226];
            n_Body_y[1226] = c_Body_y[1226];
            n_Body_x[1227] = c_Body_x[1227];
            n_Body_y[1227] = c_Body_y[1227];
            n_Body_x[1228] = c_Body_x[1228];
            n_Body_y[1228] = c_Body_y[1228];
            n_Body_x[1229] = c_Body_x[1229];
            n_Body_y[1229] = c_Body_y[1229];
            n_Body_x[1230] = c_Body_x[1230];
            n_Body_y[1230] = c_Body_y[1230];
            n_Body_x[1231] = c_Body_x[1231];
            n_Body_y[1231] = c_Body_y[1231];
            n_Body_x[1232] = c_Body_x[1232];
            n_Body_y[1232] = c_Body_y[1232];
            n_Body_x[1233] = c_Body_x[1233];
            n_Body_y[1233] = c_Body_y[1233];
            n_Body_x[1234] = c_Body_x[1234];
            n_Body_y[1234] = c_Body_y[1234];
            n_Body_x[1235] = c_Body_x[1235];
            n_Body_y[1235] = c_Body_y[1235];
            n_Body_x[1236] = c_Body_x[1236];
            n_Body_y[1236] = c_Body_y[1236];
            n_Body_x[1237] = c_Body_x[1237];
            n_Body_y[1237] = c_Body_y[1237];
            n_Body_x[1238] = c_Body_x[1238];
            n_Body_y[1238] = c_Body_y[1238];
            n_Body_x[1239] = c_Body_x[1239];
            n_Body_y[1239] = c_Body_y[1239];
            n_Body_x[1240] = c_Body_x[1240];
            n_Body_y[1240] = c_Body_y[1240];
            n_Body_x[1241] = c_Body_x[1241];
            n_Body_y[1241] = c_Body_y[1241];
            n_Body_x[1242] = c_Body_x[1242];
            n_Body_y[1242] = c_Body_y[1242];
            n_Body_x[1243] = c_Body_x[1243];
            n_Body_y[1243] = c_Body_y[1243];
            n_Body_x[1244] = c_Body_x[1244];
            n_Body_y[1244] = c_Body_y[1244];
            n_Body_x[1245] = c_Body_x[1245];
            n_Body_y[1245] = c_Body_y[1245];
            n_Body_x[1246] = c_Body_x[1246];
            n_Body_y[1246] = c_Body_y[1246];
            n_Body_x[1247] = c_Body_x[1247];
            n_Body_y[1247] = c_Body_y[1247];
            n_Body_x[1248] = c_Body_x[1248];
            n_Body_y[1248] = c_Body_y[1248];
            n_Body_x[1249] = c_Body_x[1249];
            n_Body_y[1249] = c_Body_y[1249];
            n_Body_x[1250] = c_Body_x[1250];
            n_Body_y[1250] = c_Body_y[1250];
            n_Body_x[1251] = c_Body_x[1251];
            n_Body_y[1251] = c_Body_y[1251];
            n_Body_x[1252] = c_Body_x[1252];
            n_Body_y[1252] = c_Body_y[1252];
            n_Body_x[1253] = c_Body_x[1253];
            n_Body_y[1253] = c_Body_y[1253];
            n_Body_x[1254] = c_Body_x[1254];
            n_Body_y[1254] = c_Body_y[1254];
            n_Body_x[1255] = c_Body_x[1255];
            n_Body_y[1255] = c_Body_y[1255];
            n_Body_x[1256] = c_Body_x[1256];
            n_Body_y[1256] = c_Body_y[1256];
            n_Body_x[1257] = c_Body_x[1257];
            n_Body_y[1257] = c_Body_y[1257];
            n_Body_x[1258] = c_Body_x[1258];
            n_Body_y[1258] = c_Body_y[1258];
            n_Body_x[1259] = c_Body_x[1259];
            n_Body_y[1259] = c_Body_y[1259];
            n_Body_x[1260] = c_Body_x[1260];
            n_Body_y[1260] = c_Body_y[1260];
            n_Body_x[1261] = c_Body_x[1261];
            n_Body_y[1261] = c_Body_y[1261];
            n_Body_x[1262] = c_Body_x[1262];
            n_Body_y[1262] = c_Body_y[1262];
            n_Body_x[1263] = c_Body_x[1263];
            n_Body_y[1263] = c_Body_y[1263];
            n_Body_x[1264] = c_Body_x[1264];
            n_Body_y[1264] = c_Body_y[1264];
            n_Body_x[1265] = c_Body_x[1265];
            n_Body_y[1265] = c_Body_y[1265];
            n_Body_x[1266] = c_Body_x[1266];
            n_Body_y[1266] = c_Body_y[1266];
            n_Body_x[1267] = c_Body_x[1267];
            n_Body_y[1267] = c_Body_y[1267];
            n_Body_x[1268] = c_Body_x[1268];
            n_Body_y[1268] = c_Body_y[1268];
            n_Body_x[1269] = c_Body_x[1269];
            n_Body_y[1269] = c_Body_y[1269];
            n_Body_x[1270] = c_Body_x[1270];
            n_Body_y[1270] = c_Body_y[1270];
            n_Body_x[1271] = c_Body_x[1271];
            n_Body_y[1271] = c_Body_y[1271];
            n_Body_x[1272] = c_Body_x[1272];
            n_Body_y[1272] = c_Body_y[1272];
            n_Body_x[1273] = c_Body_x[1273];
            n_Body_y[1273] = c_Body_y[1273];
            n_Body_x[1274] = c_Body_x[1274];
            n_Body_y[1274] = c_Body_y[1274];
            n_Body_x[1275] = c_Body_x[1275];
            n_Body_y[1275] = c_Body_y[1275];
            n_Body_x[1276] = c_Body_x[1276];
            n_Body_y[1276] = c_Body_y[1276];
            n_Body_x[1277] = c_Body_x[1277];
            n_Body_y[1277] = c_Body_y[1277];
            n_Body_x[1278] = c_Body_x[1278];
            n_Body_y[1278] = c_Body_y[1278];
            n_Body_x[1279] = c_Body_x[1279];
            n_Body_y[1279] = c_Body_y[1279];
            n_Body_x[1280] = c_Body_x[1280];
            n_Body_y[1280] = c_Body_y[1280];
            n_Body_x[1281] = c_Body_x[1281];
            n_Body_y[1281] = c_Body_y[1281];
            n_Body_x[1282] = c_Body_x[1282];
            n_Body_y[1282] = c_Body_y[1282];
            n_Body_x[1283] = c_Body_x[1283];
            n_Body_y[1283] = c_Body_y[1283];
            n_Body_x[1284] = c_Body_x[1284];
            n_Body_y[1284] = c_Body_y[1284];
            n_Body_x[1285] = c_Body_x[1285];
            n_Body_y[1285] = c_Body_y[1285];
            n_Body_x[1286] = c_Body_x[1286];
            n_Body_y[1286] = c_Body_y[1286];
            n_Body_x[1287] = c_Body_x[1287];
            n_Body_y[1287] = c_Body_y[1287];
            n_Body_x[1288] = c_Body_x[1288];
            n_Body_y[1288] = c_Body_y[1288];
            n_Body_x[1289] = c_Body_x[1289];
            n_Body_y[1289] = c_Body_y[1289];
            n_Body_x[1290] = c_Body_x[1290];
            n_Body_y[1290] = c_Body_y[1290];
            n_Body_x[1291] = c_Body_x[1291];
            n_Body_y[1291] = c_Body_y[1291];
            n_Body_x[1292] = c_Body_x[1292];
            n_Body_y[1292] = c_Body_y[1292];
            n_Body_x[1293] = c_Body_x[1293];
            n_Body_y[1293] = c_Body_y[1293];
            n_Body_x[1294] = c_Body_x[1294];
            n_Body_y[1294] = c_Body_y[1294];
            n_Body_x[1295] = c_Body_x[1295];
            n_Body_y[1295] = c_Body_y[1295];
            n_Body_x[1296] = c_Body_x[1296];
            n_Body_y[1296] = c_Body_y[1296];
            n_Body_x[1297] = c_Body_x[1297];
            n_Body_y[1297] = c_Body_y[1297];
            n_Body_x[1298] = c_Body_x[1298];
            n_Body_y[1298] = c_Body_y[1298];
            n_Body_x[1299] = c_Body_x[1299];
            n_Body_y[1299] = c_Body_y[1299];
            n_Body_x[1300] = c_Body_x[1300];
            n_Body_y[1300] = c_Body_y[1300];
            n_Body_x[1301] = c_Body_x[1301];
            n_Body_y[1301] = c_Body_y[1301];
            n_Body_x[1302] = c_Body_x[1302];
            n_Body_y[1302] = c_Body_y[1302];
            n_Body_x[1303] = c_Body_x[1303];
            n_Body_y[1303] = c_Body_y[1303];
            n_Body_x[1304] = c_Body_x[1304];
            n_Body_y[1304] = c_Body_y[1304];
            n_Body_x[1305] = c_Body_x[1305];
            n_Body_y[1305] = c_Body_y[1305];
            n_Body_x[1306] = c_Body_x[1306];
            n_Body_y[1306] = c_Body_y[1306];
            n_Body_x[1307] = c_Body_x[1307];
            n_Body_y[1307] = c_Body_y[1307];
            n_Body_x[1308] = c_Body_x[1308];
            n_Body_y[1308] = c_Body_y[1308];
            n_Body_x[1309] = c_Body_x[1309];
            n_Body_y[1309] = c_Body_y[1309];
            n_Body_x[1310] = c_Body_x[1310];
            n_Body_y[1310] = c_Body_y[1310];
            n_Body_x[1311] = c_Body_x[1311];
            n_Body_y[1311] = c_Body_y[1311];
            n_Body_x[1312] = c_Body_x[1312];
            n_Body_y[1312] = c_Body_y[1312];
            n_Body_x[1313] = c_Body_x[1313];
            n_Body_y[1313] = c_Body_y[1313];
            n_Body_x[1314] = c_Body_x[1314];
            n_Body_y[1314] = c_Body_y[1314];
            n_Body_x[1315] = c_Body_x[1315];
            n_Body_y[1315] = c_Body_y[1315];
            n_Body_x[1316] = c_Body_x[1316];
            n_Body_y[1316] = c_Body_y[1316];
            n_Body_x[1317] = c_Body_x[1317];
            n_Body_y[1317] = c_Body_y[1317];
            n_Body_x[1318] = c_Body_x[1318];
            n_Body_y[1318] = c_Body_y[1318];
            n_Body_x[1319] = c_Body_x[1319];
            n_Body_y[1319] = c_Body_y[1319];
            n_Body_x[1320] = c_Body_x[1320];
            n_Body_y[1320] = c_Body_y[1320];
            n_Body_x[1321] = c_Body_x[1321];
            n_Body_y[1321] = c_Body_y[1321];
            n_Body_x[1322] = c_Body_x[1322];
            n_Body_y[1322] = c_Body_y[1322];
            n_Body_x[1323] = c_Body_x[1323];
            n_Body_y[1323] = c_Body_y[1323];
            n_Body_x[1324] = c_Body_x[1324];
            n_Body_y[1324] = c_Body_y[1324];
            n_Body_x[1325] = c_Body_x[1325];
            n_Body_y[1325] = c_Body_y[1325];
            n_Body_x[1326] = c_Body_x[1326];
            n_Body_y[1326] = c_Body_y[1326];
            n_Body_x[1327] = c_Body_x[1327];
            n_Body_y[1327] = c_Body_y[1327];
            n_Body_x[1328] = c_Body_x[1328];
            n_Body_y[1328] = c_Body_y[1328];
            n_Body_x[1329] = c_Body_x[1329];
            n_Body_y[1329] = c_Body_y[1329];
            n_Body_x[1330] = c_Body_x[1330];
            n_Body_y[1330] = c_Body_y[1330];
            n_Body_x[1331] = c_Body_x[1331];
            n_Body_y[1331] = c_Body_y[1331];
            n_Body_x[1332] = c_Body_x[1332];
            n_Body_y[1332] = c_Body_y[1332];
            n_Body_x[1333] = c_Body_x[1333];
            n_Body_y[1333] = c_Body_y[1333];
            n_Body_x[1334] = c_Body_x[1334];
            n_Body_y[1334] = c_Body_y[1334];
            n_Body_x[1335] = c_Body_x[1335];
            n_Body_y[1335] = c_Body_y[1335];
            n_Body_x[1336] = c_Body_x[1336];
            n_Body_y[1336] = c_Body_y[1336];
            n_Body_x[1337] = c_Body_x[1337];
            n_Body_y[1337] = c_Body_y[1337];
            n_Body_x[1338] = c_Body_x[1338];
            n_Body_y[1338] = c_Body_y[1338];
            n_Body_x[1339] = c_Body_x[1339];
            n_Body_y[1339] = c_Body_y[1339];
            n_Body_x[1340] = c_Body_x[1340];
            n_Body_y[1340] = c_Body_y[1340];
            n_Body_x[1341] = c_Body_x[1341];
            n_Body_y[1341] = c_Body_y[1341];
            n_Body_x[1342] = c_Body_x[1342];
            n_Body_y[1342] = c_Body_y[1342];
            n_Body_x[1343] = c_Body_x[1343];
            n_Body_y[1343] = c_Body_y[1343];
            n_Body_x[1344] = c_Body_x[1344];
            n_Body_y[1344] = c_Body_y[1344];
            n_Body_x[1345] = c_Body_x[1345];
            n_Body_y[1345] = c_Body_y[1345];
            n_Body_x[1346] = c_Body_x[1346];
            n_Body_y[1346] = c_Body_y[1346];
            n_Body_x[1347] = c_Body_x[1347];
            n_Body_y[1347] = c_Body_y[1347];
            n_Body_x[1348] = c_Body_x[1348];
            n_Body_y[1348] = c_Body_y[1348];
            n_Body_x[1349] = c_Body_x[1349];
            n_Body_y[1349] = c_Body_y[1349];
            n_Body_x[1350] = c_Body_x[1350];
            n_Body_y[1350] = c_Body_y[1350];
            n_Body_x[1351] = c_Body_x[1351];
            n_Body_y[1351] = c_Body_y[1351];
            n_Body_x[1352] = c_Body_x[1352];
            n_Body_y[1352] = c_Body_y[1352];
            n_Body_x[1353] = c_Body_x[1353];
            n_Body_y[1353] = c_Body_y[1353];
            n_Body_x[1354] = c_Body_x[1354];
            n_Body_y[1354] = c_Body_y[1354];
            n_Body_x[1355] = c_Body_x[1355];
            n_Body_y[1355] = c_Body_y[1355];
            n_Body_x[1356] = c_Body_x[1356];
            n_Body_y[1356] = c_Body_y[1356];
            n_Body_x[1357] = c_Body_x[1357];
            n_Body_y[1357] = c_Body_y[1357];
            n_Body_x[1358] = c_Body_x[1358];
            n_Body_y[1358] = c_Body_y[1358];
            n_Body_x[1359] = c_Body_x[1359];
            n_Body_y[1359] = c_Body_y[1359];
            n_Body_x[1360] = c_Body_x[1360];
            n_Body_y[1360] = c_Body_y[1360];
            n_Body_x[1361] = c_Body_x[1361];
            n_Body_y[1361] = c_Body_y[1361];
            n_Body_x[1362] = c_Body_x[1362];
            n_Body_y[1362] = c_Body_y[1362];
            n_Body_x[1363] = c_Body_x[1363];
            n_Body_y[1363] = c_Body_y[1363];
            n_Body_x[1364] = c_Body_x[1364];
            n_Body_y[1364] = c_Body_y[1364];
            n_Body_x[1365] = c_Body_x[1365];
            n_Body_y[1365] = c_Body_y[1365];
            n_Body_x[1366] = c_Body_x[1366];
            n_Body_y[1366] = c_Body_y[1366];
            n_Body_x[1367] = c_Body_x[1367];
            n_Body_y[1367] = c_Body_y[1367];
            n_Body_x[1368] = c_Body_x[1368];
            n_Body_y[1368] = c_Body_y[1368];
            n_Body_x[1369] = c_Body_x[1369];
            n_Body_y[1369] = c_Body_y[1369];
            n_Body_x[1370] = c_Body_x[1370];
            n_Body_y[1370] = c_Body_y[1370];
            n_Body_x[1371] = c_Body_x[1371];
            n_Body_y[1371] = c_Body_y[1371];
            n_Body_x[1372] = c_Body_x[1372];
            n_Body_y[1372] = c_Body_y[1372];
            n_Body_x[1373] = c_Body_x[1373];
            n_Body_y[1373] = c_Body_y[1373];
            n_Body_x[1374] = c_Body_x[1374];
            n_Body_y[1374] = c_Body_y[1374];
            n_Body_x[1375] = c_Body_x[1375];
            n_Body_y[1375] = c_Body_y[1375];
            n_Body_x[1376] = c_Body_x[1376];
            n_Body_y[1376] = c_Body_y[1376];
            n_Body_x[1377] = c_Body_x[1377];
            n_Body_y[1377] = c_Body_y[1377];
            n_Body_x[1378] = c_Body_x[1378];
            n_Body_y[1378] = c_Body_y[1378];
            n_Body_x[1379] = c_Body_x[1379];
            n_Body_y[1379] = c_Body_y[1379];
            n_Body_x[1380] = c_Body_x[1380];
            n_Body_y[1380] = c_Body_y[1380];
            n_Body_x[1381] = c_Body_x[1381];
            n_Body_y[1381] = c_Body_y[1381];
            n_Body_x[1382] = c_Body_x[1382];
            n_Body_y[1382] = c_Body_y[1382];
            n_Body_x[1383] = c_Body_x[1383];
            n_Body_y[1383] = c_Body_y[1383];
            n_Body_x[1384] = c_Body_x[1384];
            n_Body_y[1384] = c_Body_y[1384];
            n_Body_x[1385] = c_Body_x[1385];
            n_Body_y[1385] = c_Body_y[1385];
            n_Body_x[1386] = c_Body_x[1386];
            n_Body_y[1386] = c_Body_y[1386];
            n_Body_x[1387] = c_Body_x[1387];
            n_Body_y[1387] = c_Body_y[1387];
            n_Body_x[1388] = c_Body_x[1388];
            n_Body_y[1388] = c_Body_y[1388];
            n_Body_x[1389] = c_Body_x[1389];
            n_Body_y[1389] = c_Body_y[1389];
            n_Body_x[1390] = c_Body_x[1390];
            n_Body_y[1390] = c_Body_y[1390];
            n_Body_x[1391] = c_Body_x[1391];
            n_Body_y[1391] = c_Body_y[1391];
            n_Body_x[1392] = c_Body_x[1392];
            n_Body_y[1392] = c_Body_y[1392];
            n_Body_x[1393] = c_Body_x[1393];
            n_Body_y[1393] = c_Body_y[1393];
            n_Body_x[1394] = c_Body_x[1394];
            n_Body_y[1394] = c_Body_y[1394];
            n_Body_x[1395] = c_Body_x[1395];
            n_Body_y[1395] = c_Body_y[1395];
            n_Body_x[1396] = c_Body_x[1396];
            n_Body_y[1396] = c_Body_y[1396];
            n_Body_x[1397] = c_Body_x[1397];
            n_Body_y[1397] = c_Body_y[1397];
            n_Body_x[1398] = c_Body_x[1398];
            n_Body_y[1398] = c_Body_y[1398];
            n_Body_x[1399] = c_Body_x[1399];
            n_Body_y[1399] = c_Body_y[1399];
            n_Body_x[1400] = c_Body_x[1400];
            n_Body_y[1400] = c_Body_y[1400];
            n_Body_x[1401] = c_Body_x[1401];
            n_Body_y[1401] = c_Body_y[1401];
            n_Body_x[1402] = c_Body_x[1402];
            n_Body_y[1402] = c_Body_y[1402];
            n_Body_x[1403] = c_Body_x[1403];
            n_Body_y[1403] = c_Body_y[1403];
            n_Body_x[1404] = c_Body_x[1404];
            n_Body_y[1404] = c_Body_y[1404];
            n_Body_x[1405] = c_Body_x[1405];
            n_Body_y[1405] = c_Body_y[1405];
            n_Body_x[1406] = c_Body_x[1406];
            n_Body_y[1406] = c_Body_y[1406];
            n_Body_x[1407] = c_Body_x[1407];
            n_Body_y[1407] = c_Body_y[1407];
            n_Body_x[1408] = c_Body_x[1408];
            n_Body_y[1408] = c_Body_y[1408];
            n_Body_x[1409] = c_Body_x[1409];
            n_Body_y[1409] = c_Body_y[1409];
            n_Body_x[1410] = c_Body_x[1410];
            n_Body_y[1410] = c_Body_y[1410];
            n_Body_x[1411] = c_Body_x[1411];
            n_Body_y[1411] = c_Body_y[1411];
            n_Body_x[1412] = c_Body_x[1412];
            n_Body_y[1412] = c_Body_y[1412];
            n_Body_x[1413] = c_Body_x[1413];
            n_Body_y[1413] = c_Body_y[1413];
            n_Body_x[1414] = c_Body_x[1414];
            n_Body_y[1414] = c_Body_y[1414];
            n_Body_x[1415] = c_Body_x[1415];
            n_Body_y[1415] = c_Body_y[1415];
            n_Body_x[1416] = c_Body_x[1416];
            n_Body_y[1416] = c_Body_y[1416];
            n_Body_x[1417] = c_Body_x[1417];
            n_Body_y[1417] = c_Body_y[1417];
            n_Body_x[1418] = c_Body_x[1418];
            n_Body_y[1418] = c_Body_y[1418];
            n_Body_x[1419] = c_Body_x[1419];
            n_Body_y[1419] = c_Body_y[1419];
            n_Body_x[1420] = c_Body_x[1420];
            n_Body_y[1420] = c_Body_y[1420];
            n_Body_x[1421] = c_Body_x[1421];
            n_Body_y[1421] = c_Body_y[1421];
            n_Body_x[1422] = c_Body_x[1422];
            n_Body_y[1422] = c_Body_y[1422];
            n_Body_x[1423] = c_Body_x[1423];
            n_Body_y[1423] = c_Body_y[1423];
            n_Body_x[1424] = c_Body_x[1424];
            n_Body_y[1424] = c_Body_y[1424];
            n_Body_x[1425] = c_Body_x[1425];
            n_Body_y[1425] = c_Body_y[1425];
            n_Body_x[1426] = c_Body_x[1426];
            n_Body_y[1426] = c_Body_y[1426];
            n_Body_x[1427] = c_Body_x[1427];
            n_Body_y[1427] = c_Body_y[1427];
            n_Body_x[1428] = c_Body_x[1428];
            n_Body_y[1428] = c_Body_y[1428];
            n_Body_x[1429] = c_Body_x[1429];
            n_Body_y[1429] = c_Body_y[1429];
            n_Body_x[1430] = c_Body_x[1430];
            n_Body_y[1430] = c_Body_y[1430];
            n_Body_x[1431] = c_Body_x[1431];
            n_Body_y[1431] = c_Body_y[1431];
            n_Body_x[1432] = c_Body_x[1432];
            n_Body_y[1432] = c_Body_y[1432];
            n_Body_x[1433] = c_Body_x[1433];
            n_Body_y[1433] = c_Body_y[1433];
            n_Body_x[1434] = c_Body_x[1434];
            n_Body_y[1434] = c_Body_y[1434];
            n_Body_x[1435] = c_Body_x[1435];
            n_Body_y[1435] = c_Body_y[1435];
            n_Body_x[1436] = c_Body_x[1436];
            n_Body_y[1436] = c_Body_y[1436];
            n_Body_x[1437] = c_Body_x[1437];
            n_Body_y[1437] = c_Body_y[1437];
            n_Body_x[1438] = c_Body_x[1438];
            n_Body_y[1438] = c_Body_y[1438];
            n_Body_x[1439] = c_Body_x[1439];
            n_Body_y[1439] = c_Body_y[1439];
            n_Body_x[1440] = c_Body_x[1440];
            n_Body_y[1440] = c_Body_y[1440];
            n_Body_x[1441] = c_Body_x[1441];
            n_Body_y[1441] = c_Body_y[1441];
            n_Body_x[1442] = c_Body_x[1442];
            n_Body_y[1442] = c_Body_y[1442];
            n_Body_x[1443] = c_Body_x[1443];
            n_Body_y[1443] = c_Body_y[1443];
            n_Body_x[1444] = c_Body_x[1444];
            n_Body_y[1444] = c_Body_y[1444];
            n_Body_x[1445] = c_Body_x[1445];
            n_Body_y[1445] = c_Body_y[1445];
            n_Body_x[1446] = c_Body_x[1446];
            n_Body_y[1446] = c_Body_y[1446];
            n_Body_x[1447] = c_Body_x[1447];
            n_Body_y[1447] = c_Body_y[1447];
            n_Body_x[1448] = c_Body_x[1448];
            n_Body_y[1448] = c_Body_y[1448];
            n_Body_x[1449] = c_Body_x[1449];
            n_Body_y[1449] = c_Body_y[1449];
            n_Body_x[1450] = c_Body_x[1450];
            n_Body_y[1450] = c_Body_y[1450];
            n_Body_x[1451] = c_Body_x[1451];
            n_Body_y[1451] = c_Body_y[1451];
            n_Body_x[1452] = c_Body_x[1452];
            n_Body_y[1452] = c_Body_y[1452];
            n_Body_x[1453] = c_Body_x[1453];
            n_Body_y[1453] = c_Body_y[1453];
            n_Body_x[1454] = c_Body_x[1454];
            n_Body_y[1454] = c_Body_y[1454];
            n_Body_x[1455] = c_Body_x[1455];
            n_Body_y[1455] = c_Body_y[1455];
            n_Body_x[1456] = c_Body_x[1456];
            n_Body_y[1456] = c_Body_y[1456];
            n_Body_x[1457] = c_Body_x[1457];
            n_Body_y[1457] = c_Body_y[1457];
            n_Body_x[1458] = c_Body_x[1458];
            n_Body_y[1458] = c_Body_y[1458];
            n_Body_x[1459] = c_Body_x[1459];
            n_Body_y[1459] = c_Body_y[1459];
            n_Body_x[1460] = c_Body_x[1460];
            n_Body_y[1460] = c_Body_y[1460];
            n_Body_x[1461] = c_Body_x[1461];
            n_Body_y[1461] = c_Body_y[1461];
            n_Body_x[1462] = c_Body_x[1462];
            n_Body_y[1462] = c_Body_y[1462];
            n_Body_x[1463] = c_Body_x[1463];
            n_Body_y[1463] = c_Body_y[1463];
            n_Body_x[1464] = c_Body_x[1464];
            n_Body_y[1464] = c_Body_y[1464];
            n_Body_x[1465] = c_Body_x[1465];
            n_Body_y[1465] = c_Body_y[1465];
            n_Body_x[1466] = c_Body_x[1466];
            n_Body_y[1466] = c_Body_y[1466];
            n_Body_x[1467] = c_Body_x[1467];
            n_Body_y[1467] = c_Body_y[1467];
            n_Body_x[1468] = c_Body_x[1468];
            n_Body_y[1468] = c_Body_y[1468];
            n_Body_x[1469] = c_Body_x[1469];
            n_Body_y[1469] = c_Body_y[1469];
            n_Body_x[1470] = c_Body_x[1470];
            n_Body_y[1470] = c_Body_y[1470];
            n_Body_x[1471] = c_Body_x[1471];
            n_Body_y[1471] = c_Body_y[1471];
            n_Body_x[1472] = c_Body_x[1472];
            n_Body_y[1472] = c_Body_y[1472];
            n_Body_x[1473] = c_Body_x[1473];
            n_Body_y[1473] = c_Body_y[1473];
            n_Body_x[1474] = c_Body_x[1474];
            n_Body_y[1474] = c_Body_y[1474];
            n_Body_x[1475] = c_Body_x[1475];
            n_Body_y[1475] = c_Body_y[1475];
            n_Body_x[1476] = c_Body_x[1476];
            n_Body_y[1476] = c_Body_y[1476];
            n_Body_x[1477] = c_Body_x[1477];
            n_Body_y[1477] = c_Body_y[1477];
            n_Body_x[1478] = c_Body_x[1478];
            n_Body_y[1478] = c_Body_y[1478];
            n_Body_x[1479] = c_Body_x[1479];
            n_Body_y[1479] = c_Body_y[1479];
            n_Body_x[1480] = c_Body_x[1480];
            n_Body_y[1480] = c_Body_y[1480];
            n_Body_x[1481] = c_Body_x[1481];
            n_Body_y[1481] = c_Body_y[1481];
            n_Body_x[1482] = c_Body_x[1482];
            n_Body_y[1482] = c_Body_y[1482];
            n_Body_x[1483] = c_Body_x[1483];
            n_Body_y[1483] = c_Body_y[1483];
            n_Body_x[1484] = c_Body_x[1484];
            n_Body_y[1484] = c_Body_y[1484];
            n_Body_x[1485] = c_Body_x[1485];
            n_Body_y[1485] = c_Body_y[1485];
            n_Body_x[1486] = c_Body_x[1486];
            n_Body_y[1486] = c_Body_y[1486];
            n_Body_x[1487] = c_Body_x[1487];
            n_Body_y[1487] = c_Body_y[1487];
            n_Body_x[1488] = c_Body_x[1488];
            n_Body_y[1488] = c_Body_y[1488];
            n_Body_x[1489] = c_Body_x[1489];
            n_Body_y[1489] = c_Body_y[1489];
            n_Body_x[1490] = c_Body_x[1490];
            n_Body_y[1490] = c_Body_y[1490];
            n_Body_x[1491] = c_Body_x[1491];
            n_Body_y[1491] = c_Body_y[1491];
            n_Body_x[1492] = c_Body_x[1492];
            n_Body_y[1492] = c_Body_y[1492];
            n_Body_x[1493] = c_Body_x[1493];
            n_Body_y[1493] = c_Body_y[1493];
            n_Body_x[1494] = c_Body_x[1494];
            n_Body_y[1494] = c_Body_y[1494];
            n_Body_x[1495] = c_Body_x[1495];
            n_Body_y[1495] = c_Body_y[1495];
            n_Body_x[1496] = c_Body_x[1496];
            n_Body_y[1496] = c_Body_y[1496];
            n_Body_x[1497] = c_Body_x[1497];
            n_Body_y[1497] = c_Body_y[1497];
            n_Body_x[1498] = c_Body_x[1498];
            n_Body_y[1498] = c_Body_y[1498];
            n_Body_x[1499] = c_Body_x[1499];
            n_Body_y[1499] = c_Body_y[1499];
            n_Body_x[1500] = c_Body_x[1500];
            n_Body_y[1500] = c_Body_y[1500];
            n_Body_x[1501] = c_Body_x[1501];
            n_Body_y[1501] = c_Body_y[1501];
            n_Body_x[1502] = c_Body_x[1502];
            n_Body_y[1502] = c_Body_y[1502];
            n_Body_x[1503] = c_Body_x[1503];
            n_Body_y[1503] = c_Body_y[1503];
            n_Body_x[1504] = c_Body_x[1504];
            n_Body_y[1504] = c_Body_y[1504];
            n_Body_x[1505] = c_Body_x[1505];
            n_Body_y[1505] = c_Body_y[1505];
            n_Body_x[1506] = c_Body_x[1506];
            n_Body_y[1506] = c_Body_y[1506];
            n_Body_x[1507] = c_Body_x[1507];
            n_Body_y[1507] = c_Body_y[1507];
            n_Body_x[1508] = c_Body_x[1508];
            n_Body_y[1508] = c_Body_y[1508];
            n_Body_x[1509] = c_Body_x[1509];
            n_Body_y[1509] = c_Body_y[1509];
            n_Body_x[1510] = c_Body_x[1510];
            n_Body_y[1510] = c_Body_y[1510];
            n_Body_x[1511] = c_Body_x[1511];
            n_Body_y[1511] = c_Body_y[1511];
            n_Body_x[1512] = c_Body_x[1512];
            n_Body_y[1512] = c_Body_y[1512];
            n_Body_x[1513] = c_Body_x[1513];
            n_Body_y[1513] = c_Body_y[1513];
            n_Body_x[1514] = c_Body_x[1514];
            n_Body_y[1514] = c_Body_y[1514];
            n_Body_x[1515] = c_Body_x[1515];
            n_Body_y[1515] = c_Body_y[1515];
            n_Body_x[1516] = c_Body_x[1516];
            n_Body_y[1516] = c_Body_y[1516];
            n_Body_x[1517] = c_Body_x[1517];
            n_Body_y[1517] = c_Body_y[1517];
            n_Body_x[1518] = c_Body_x[1518];
            n_Body_y[1518] = c_Body_y[1518];
            n_Body_x[1519] = c_Body_x[1519];
            n_Body_y[1519] = c_Body_y[1519];
            n_Body_x[1520] = c_Body_x[1520];
            n_Body_y[1520] = c_Body_y[1520];
            n_Body_x[1521] = c_Body_x[1521];
            n_Body_y[1521] = c_Body_y[1521];
            n_Body_x[1522] = c_Body_x[1522];
            n_Body_y[1522] = c_Body_y[1522];
            n_Body_x[1523] = c_Body_x[1523];
            n_Body_y[1523] = c_Body_y[1523];
            n_Body_x[1524] = c_Body_x[1524];
            n_Body_y[1524] = c_Body_y[1524];
            n_Body_x[1525] = c_Body_x[1525];
            n_Body_y[1525] = c_Body_y[1525];
            n_Body_x[1526] = c_Body_x[1526];
            n_Body_y[1526] = c_Body_y[1526];
            n_Body_x[1527] = c_Body_x[1527];
            n_Body_y[1527] = c_Body_y[1527];
            n_Body_x[1528] = c_Body_x[1528];
            n_Body_y[1528] = c_Body_y[1528];
            n_Body_x[1529] = c_Body_x[1529];
            n_Body_y[1529] = c_Body_y[1529];
            n_Body_x[1530] = c_Body_x[1530];
            n_Body_y[1530] = c_Body_y[1530];
            n_Body_x[1531] = c_Body_x[1531];
            n_Body_y[1531] = c_Body_y[1531];
            n_Body_x[1532] = c_Body_x[1532];
            n_Body_y[1532] = c_Body_y[1532];
            n_Body_x[1533] = c_Body_x[1533];
            n_Body_y[1533] = c_Body_y[1533];
            n_Body_x[1534] = c_Body_x[1534];
            n_Body_y[1534] = c_Body_y[1534];
            n_Body_x[1535] = c_Body_x[1535];
            n_Body_y[1535] = c_Body_y[1535];
            n_Body_x[1536] = c_Body_x[1536];
            n_Body_y[1536] = c_Body_y[1536];
            n_Body_x[1537] = c_Body_x[1537];
            n_Body_y[1537] = c_Body_y[1537];
            n_Body_x[1538] = c_Body_x[1538];
            n_Body_y[1538] = c_Body_y[1538];
            n_Body_x[1539] = c_Body_x[1539];
            n_Body_y[1539] = c_Body_y[1539];
            n_Body_x[1540] = c_Body_x[1540];
            n_Body_y[1540] = c_Body_y[1540];
            n_Body_x[1541] = c_Body_x[1541];
            n_Body_y[1541] = c_Body_y[1541];
            n_Body_x[1542] = c_Body_x[1542];
            n_Body_y[1542] = c_Body_y[1542];
            n_Body_x[1543] = c_Body_x[1543];
            n_Body_y[1543] = c_Body_y[1543];
            n_Body_x[1544] = c_Body_x[1544];
            n_Body_y[1544] = c_Body_y[1544];
            n_Body_x[1545] = c_Body_x[1545];
            n_Body_y[1545] = c_Body_y[1545];
            n_Body_x[1546] = c_Body_x[1546];
            n_Body_y[1546] = c_Body_y[1546];
            n_Body_x[1547] = c_Body_x[1547];
            n_Body_y[1547] = c_Body_y[1547];
            n_Body_x[1548] = c_Body_x[1548];
            n_Body_y[1548] = c_Body_y[1548];
            n_Body_x[1549] = c_Body_x[1549];
            n_Body_y[1549] = c_Body_y[1549];
            n_Body_x[1550] = c_Body_x[1550];
            n_Body_y[1550] = c_Body_y[1550];
            n_Body_x[1551] = c_Body_x[1551];
            n_Body_y[1551] = c_Body_y[1551];
            n_Body_x[1552] = c_Body_x[1552];
            n_Body_y[1552] = c_Body_y[1552];
            n_Body_x[1553] = c_Body_x[1553];
            n_Body_y[1553] = c_Body_y[1553];
            n_Body_x[1554] = c_Body_x[1554];
            n_Body_y[1554] = c_Body_y[1554];
            n_Body_x[1555] = c_Body_x[1555];
            n_Body_y[1555] = c_Body_y[1555];
            n_Body_x[1556] = c_Body_x[1556];
            n_Body_y[1556] = c_Body_y[1556];
            n_Body_x[1557] = c_Body_x[1557];
            n_Body_y[1557] = c_Body_y[1557];
            n_Body_x[1558] = c_Body_x[1558];
            n_Body_y[1558] = c_Body_y[1558];
            n_Body_x[1559] = c_Body_x[1559];
            n_Body_y[1559] = c_Body_y[1559];
            n_Body_x[1560] = c_Body_x[1560];
            n_Body_y[1560] = c_Body_y[1560];
            n_Body_x[1561] = c_Body_x[1561];
            n_Body_y[1561] = c_Body_y[1561];
            n_Body_x[1562] = c_Body_x[1562];
            n_Body_y[1562] = c_Body_y[1562];
            n_Body_x[1563] = c_Body_x[1563];
            n_Body_y[1563] = c_Body_y[1563];
            n_Body_x[1564] = c_Body_x[1564];
            n_Body_y[1564] = c_Body_y[1564];
            n_Body_x[1565] = c_Body_x[1565];
            n_Body_y[1565] = c_Body_y[1565];
            n_Body_x[1566] = c_Body_x[1566];
            n_Body_y[1566] = c_Body_y[1566];
            n_Body_x[1567] = c_Body_x[1567];
            n_Body_y[1567] = c_Body_y[1567];
            n_Body_x[1568] = c_Body_x[1568];
            n_Body_y[1568] = c_Body_y[1568];
            n_Body_x[1569] = c_Body_x[1569];
            n_Body_y[1569] = c_Body_y[1569];
            n_Body_x[1570] = c_Body_x[1570];
            n_Body_y[1570] = c_Body_y[1570];
            n_Body_x[1571] = c_Body_x[1571];
            n_Body_y[1571] = c_Body_y[1571];
            n_Body_x[1572] = c_Body_x[1572];
            n_Body_y[1572] = c_Body_y[1572];
            n_Body_x[1573] = c_Body_x[1573];
            n_Body_y[1573] = c_Body_y[1573];
            n_Body_x[1574] = c_Body_x[1574];
            n_Body_y[1574] = c_Body_y[1574];
            n_Body_x[1575] = c_Body_x[1575];
            n_Body_y[1575] = c_Body_y[1575];
            n_Body_x[1576] = c_Body_x[1576];
            n_Body_y[1576] = c_Body_y[1576];
            n_Body_x[1577] = c_Body_x[1577];
            n_Body_y[1577] = c_Body_y[1577];
            n_Body_x[1578] = c_Body_x[1578];
            n_Body_y[1578] = c_Body_y[1578];
            n_Body_x[1579] = c_Body_x[1579];
            n_Body_y[1579] = c_Body_y[1579];
            n_Body_x[1580] = c_Body_x[1580];
            n_Body_y[1580] = c_Body_y[1580];
            n_Body_x[1581] = c_Body_x[1581];
            n_Body_y[1581] = c_Body_y[1581];
            n_Body_x[1582] = c_Body_x[1582];
            n_Body_y[1582] = c_Body_y[1582];
            n_Body_x[1583] = c_Body_x[1583];
            n_Body_y[1583] = c_Body_y[1583];
            n_Body_x[1584] = c_Body_x[1584];
            n_Body_y[1584] = c_Body_y[1584];
            n_Body_x[1585] = c_Body_x[1585];
            n_Body_y[1585] = c_Body_y[1585];
            n_Body_x[1586] = c_Body_x[1586];
            n_Body_y[1586] = c_Body_y[1586];
            n_Body_x[1587] = c_Body_x[1587];
            n_Body_y[1587] = c_Body_y[1587];
            n_Body_x[1588] = c_Body_x[1588];
            n_Body_y[1588] = c_Body_y[1588];
            n_Body_x[1589] = c_Body_x[1589];
            n_Body_y[1589] = c_Body_y[1589];
            n_Body_x[1590] = c_Body_x[1590];
            n_Body_y[1590] = c_Body_y[1590];
            n_Body_x[1591] = c_Body_x[1591];
            n_Body_y[1591] = c_Body_y[1591];
            n_Body_x[1592] = c_Body_x[1592];
            n_Body_y[1592] = c_Body_y[1592];
            n_Body_x[1593] = c_Body_x[1593];
            n_Body_y[1593] = c_Body_y[1593];
            n_Body_x[1594] = c_Body_x[1594];
            n_Body_y[1594] = c_Body_y[1594];
            n_Body_x[1595] = c_Body_x[1595];
            n_Body_y[1595] = c_Body_y[1595];
            n_Body_x[1596] = c_Body_x[1596];
            n_Body_y[1596] = c_Body_y[1596];
            n_Body_x[1597] = c_Body_x[1597];
            n_Body_y[1597] = c_Body_y[1597];
            n_Body_x[1598] = c_Body_x[1598];
            n_Body_y[1598] = c_Body_y[1598];
            n_Body_x[1599] = c_Body_x[1599];
            n_Body_y[1599] = c_Body_y[1599];
            n_Body_x[1600] = c_Body_x[1600];
            n_Body_y[1600] = c_Body_y[1600];
            n_Body_x[1601] = c_Body_x[1601];
            n_Body_y[1601] = c_Body_y[1601];
            n_Body_x[1602] = c_Body_x[1602];
            n_Body_y[1602] = c_Body_y[1602];
            n_Body_x[1603] = c_Body_x[1603];
            n_Body_y[1603] = c_Body_y[1603];
            n_Body_x[1604] = c_Body_x[1604];
            n_Body_y[1604] = c_Body_y[1604];
            n_Body_x[1605] = c_Body_x[1605];
            n_Body_y[1605] = c_Body_y[1605];
            n_Body_x[1606] = c_Body_x[1606];
            n_Body_y[1606] = c_Body_y[1606];
            n_Body_x[1607] = c_Body_x[1607];
            n_Body_y[1607] = c_Body_y[1607];
            n_Body_x[1608] = c_Body_x[1608];
            n_Body_y[1608] = c_Body_y[1608];
            n_Body_x[1609] = c_Body_x[1609];
            n_Body_y[1609] = c_Body_y[1609];
            n_Body_x[1610] = c_Body_x[1610];
            n_Body_y[1610] = c_Body_y[1610];
            n_Body_x[1611] = c_Body_x[1611];
            n_Body_y[1611] = c_Body_y[1611];
            n_Body_x[1612] = c_Body_x[1612];
            n_Body_y[1612] = c_Body_y[1612];
            n_Body_x[1613] = c_Body_x[1613];
            n_Body_y[1613] = c_Body_y[1613];
            n_Body_x[1614] = c_Body_x[1614];
            n_Body_y[1614] = c_Body_y[1614];
            n_Body_x[1615] = c_Body_x[1615];
            n_Body_y[1615] = c_Body_y[1615];
            n_Body_x[1616] = c_Body_x[1616];
            n_Body_y[1616] = c_Body_y[1616];
            n_Body_x[1617] = c_Body_x[1617];
            n_Body_y[1617] = c_Body_y[1617];
            n_Body_x[1618] = c_Body_x[1618];
            n_Body_y[1618] = c_Body_y[1618];
            n_Body_x[1619] = c_Body_x[1619];
            n_Body_y[1619] = c_Body_y[1619];
            n_Body_x[1620] = c_Body_x[1620];
            n_Body_y[1620] = c_Body_y[1620];
            n_Body_x[1621] = c_Body_x[1621];
            n_Body_y[1621] = c_Body_y[1621];
            n_Body_x[1622] = c_Body_x[1622];
            n_Body_y[1622] = c_Body_y[1622];
            n_Body_x[1623] = c_Body_x[1623];
            n_Body_y[1623] = c_Body_y[1623];
            n_Body_x[1624] = c_Body_x[1624];
            n_Body_y[1624] = c_Body_y[1624];
            n_Body_x[1625] = c_Body_x[1625];
            n_Body_y[1625] = c_Body_y[1625];
            n_Body_x[1626] = c_Body_x[1626];
            n_Body_y[1626] = c_Body_y[1626];
            n_Body_x[1627] = c_Body_x[1627];
            n_Body_y[1627] = c_Body_y[1627];
            n_Body_x[1628] = c_Body_x[1628];
            n_Body_y[1628] = c_Body_y[1628];
            n_Body_x[1629] = c_Body_x[1629];
            n_Body_y[1629] = c_Body_y[1629];
            n_Body_x[1630] = c_Body_x[1630];
            n_Body_y[1630] = c_Body_y[1630];
            n_Body_x[1631] = c_Body_x[1631];
            n_Body_y[1631] = c_Body_y[1631];
            n_Body_x[1632] = c_Body_x[1632];
            n_Body_y[1632] = c_Body_y[1632];
            n_Body_x[1633] = c_Body_x[1633];
            n_Body_y[1633] = c_Body_y[1633];
            n_Body_x[1634] = c_Body_x[1634];
            n_Body_y[1634] = c_Body_y[1634];
            n_Body_x[1635] = c_Body_x[1635];
            n_Body_y[1635] = c_Body_y[1635];
            n_Body_x[1636] = c_Body_x[1636];
            n_Body_y[1636] = c_Body_y[1636];
            n_Body_x[1637] = c_Body_x[1637];
            n_Body_y[1637] = c_Body_y[1637];
            n_Body_x[1638] = c_Body_x[1638];
            n_Body_y[1638] = c_Body_y[1638];
            n_Body_x[1639] = c_Body_x[1639];
            n_Body_y[1639] = c_Body_y[1639];
            n_Body_x[1640] = c_Body_x[1640];
            n_Body_y[1640] = c_Body_y[1640];
            n_Body_x[1641] = c_Body_x[1641];
            n_Body_y[1641] = c_Body_y[1641];
            n_Body_x[1642] = c_Body_x[1642];
            n_Body_y[1642] = c_Body_y[1642];
            n_Body_x[1643] = c_Body_x[1643];
            n_Body_y[1643] = c_Body_y[1643];
            n_Body_x[1644] = c_Body_x[1644];
            n_Body_y[1644] = c_Body_y[1644];
            n_Body_x[1645] = c_Body_x[1645];
            n_Body_y[1645] = c_Body_y[1645];
            n_Body_x[1646] = c_Body_x[1646];
            n_Body_y[1646] = c_Body_y[1646];
            n_Body_x[1647] = c_Body_x[1647];
            n_Body_y[1647] = c_Body_y[1647];
            n_Body_x[1648] = c_Body_x[1648];
            n_Body_y[1648] = c_Body_y[1648];
            n_Body_x[1649] = c_Body_x[1649];
            n_Body_y[1649] = c_Body_y[1649];
            n_Body_x[1650] = c_Body_x[1650];
            n_Body_y[1650] = c_Body_y[1650];
            n_Body_x[1651] = c_Body_x[1651];
            n_Body_y[1651] = c_Body_y[1651];
            n_Body_x[1652] = c_Body_x[1652];
            n_Body_y[1652] = c_Body_y[1652];
            n_Body_x[1653] = c_Body_x[1653];
            n_Body_y[1653] = c_Body_y[1653];
            n_Body_x[1654] = c_Body_x[1654];
            n_Body_y[1654] = c_Body_y[1654];
            n_Body_x[1655] = c_Body_x[1655];
            n_Body_y[1655] = c_Body_y[1655];
            n_Body_x[1656] = c_Body_x[1656];
            n_Body_y[1656] = c_Body_y[1656];
            n_Body_x[1657] = c_Body_x[1657];
            n_Body_y[1657] = c_Body_y[1657];
            n_Body_x[1658] = c_Body_x[1658];
            n_Body_y[1658] = c_Body_y[1658];
            n_Body_x[1659] = c_Body_x[1659];
            n_Body_y[1659] = c_Body_y[1659];
            n_Body_x[1660] = c_Body_x[1660];
            n_Body_y[1660] = c_Body_y[1660];
            n_Body_x[1661] = c_Body_x[1661];
            n_Body_y[1661] = c_Body_y[1661];
            n_Body_x[1662] = c_Body_x[1662];
            n_Body_y[1662] = c_Body_y[1662];
            n_Body_x[1663] = c_Body_x[1663];
            n_Body_y[1663] = c_Body_y[1663];
            n_Body_x[1664] = c_Body_x[1664];
            n_Body_y[1664] = c_Body_y[1664];
            n_Body_x[1665] = c_Body_x[1665];
            n_Body_y[1665] = c_Body_y[1665];
            n_Body_x[1666] = c_Body_x[1666];
            n_Body_y[1666] = c_Body_y[1666];
            n_Body_x[1667] = c_Body_x[1667];
            n_Body_y[1667] = c_Body_y[1667];
            n_Body_x[1668] = c_Body_x[1668];
            n_Body_y[1668] = c_Body_y[1668];
            n_Body_x[1669] = c_Body_x[1669];
            n_Body_y[1669] = c_Body_y[1669];
            n_Body_x[1670] = c_Body_x[1670];
            n_Body_y[1670] = c_Body_y[1670];
            n_Body_x[1671] = c_Body_x[1671];
            n_Body_y[1671] = c_Body_y[1671];
            n_Body_x[1672] = c_Body_x[1672];
            n_Body_y[1672] = c_Body_y[1672];
            n_Body_x[1673] = c_Body_x[1673];
            n_Body_y[1673] = c_Body_y[1673];
            n_Body_x[1674] = c_Body_x[1674];
            n_Body_y[1674] = c_Body_y[1674];
            n_Body_x[1675] = c_Body_x[1675];
            n_Body_y[1675] = c_Body_y[1675];
            n_Body_x[1676] = c_Body_x[1676];
            n_Body_y[1676] = c_Body_y[1676];
            n_Body_x[1677] = c_Body_x[1677];
            n_Body_y[1677] = c_Body_y[1677];
            n_Body_x[1678] = c_Body_x[1678];
            n_Body_y[1678] = c_Body_y[1678];
            n_Body_x[1679] = c_Body_x[1679];
            n_Body_y[1679] = c_Body_y[1679];
            n_Body_x[1680] = c_Body_x[1680];
            n_Body_y[1680] = c_Body_y[1680];
            n_Body_x[1681] = c_Body_x[1681];
            n_Body_y[1681] = c_Body_y[1681];
            n_Body_x[1682] = c_Body_x[1682];
            n_Body_y[1682] = c_Body_y[1682];
            n_Body_x[1683] = c_Body_x[1683];
            n_Body_y[1683] = c_Body_y[1683];
            n_Body_x[1684] = c_Body_x[1684];
            n_Body_y[1684] = c_Body_y[1684];
            n_Body_x[1685] = c_Body_x[1685];
            n_Body_y[1685] = c_Body_y[1685];
            n_Body_x[1686] = c_Body_x[1686];
            n_Body_y[1686] = c_Body_y[1686];
            n_Body_x[1687] = c_Body_x[1687];
            n_Body_y[1687] = c_Body_y[1687];
            n_Body_x[1688] = c_Body_x[1688];
            n_Body_y[1688] = c_Body_y[1688];
            n_Body_x[1689] = c_Body_x[1689];
            n_Body_y[1689] = c_Body_y[1689];
            n_Body_x[1690] = c_Body_x[1690];
            n_Body_y[1690] = c_Body_y[1690];
            n_Body_x[1691] = c_Body_x[1691];
            n_Body_y[1691] = c_Body_y[1691];
            n_Body_x[1692] = c_Body_x[1692];
            n_Body_y[1692] = c_Body_y[1692];
            n_Body_x[1693] = c_Body_x[1693];
            n_Body_y[1693] = c_Body_y[1693];
            n_Body_x[1694] = c_Body_x[1694];
            n_Body_y[1694] = c_Body_y[1694];
            n_Body_x[1695] = c_Body_x[1695];
            n_Body_y[1695] = c_Body_y[1695];
            n_Body_x[1696] = c_Body_x[1696];
            n_Body_y[1696] = c_Body_y[1696];
            n_Body_x[1697] = c_Body_x[1697];
            n_Body_y[1697] = c_Body_y[1697];
            n_Body_x[1698] = c_Body_x[1698];
            n_Body_y[1698] = c_Body_y[1698];
            n_Body_x[1699] = c_Body_x[1699];
            n_Body_y[1699] = c_Body_y[1699];
            n_Body_x[1700] = c_Body_x[1700];
            n_Body_y[1700] = c_Body_y[1700];
            n_Body_x[1701] = c_Body_x[1701];
            n_Body_y[1701] = c_Body_y[1701];
            n_Body_x[1702] = c_Body_x[1702];
            n_Body_y[1702] = c_Body_y[1702];
            n_Body_x[1703] = c_Body_x[1703];
            n_Body_y[1703] = c_Body_y[1703];
            n_Body_x[1704] = c_Body_x[1704];
            n_Body_y[1704] = c_Body_y[1704];
            n_Body_x[1705] = c_Body_x[1705];
            n_Body_y[1705] = c_Body_y[1705];
            n_Body_x[1706] = c_Body_x[1706];
            n_Body_y[1706] = c_Body_y[1706];
            n_Body_x[1707] = c_Body_x[1707];
            n_Body_y[1707] = c_Body_y[1707];
            n_Body_x[1708] = c_Body_x[1708];
            n_Body_y[1708] = c_Body_y[1708];
            n_Body_x[1709] = c_Body_x[1709];
            n_Body_y[1709] = c_Body_y[1709];
            n_Body_x[1710] = c_Body_x[1710];
            n_Body_y[1710] = c_Body_y[1710];
            n_Body_x[1711] = c_Body_x[1711];
            n_Body_y[1711] = c_Body_y[1711];
            n_Body_x[1712] = c_Body_x[1712];
            n_Body_y[1712] = c_Body_y[1712];
            n_Body_x[1713] = c_Body_x[1713];
            n_Body_y[1713] = c_Body_y[1713];
            n_Body_x[1714] = c_Body_x[1714];
            n_Body_y[1714] = c_Body_y[1714];
            n_Body_x[1715] = c_Body_x[1715];
            n_Body_y[1715] = c_Body_y[1715];
            n_Body_x[1716] = c_Body_x[1716];
            n_Body_y[1716] = c_Body_y[1716];
            n_Body_x[1717] = c_Body_x[1717];
            n_Body_y[1717] = c_Body_y[1717];
            n_Body_x[1718] = c_Body_x[1718];
            n_Body_y[1718] = c_Body_y[1718];
            n_Body_x[1719] = c_Body_x[1719];
            n_Body_y[1719] = c_Body_y[1719];
            n_Body_x[1720] = c_Body_x[1720];
            n_Body_y[1720] = c_Body_y[1720];
            n_Body_x[1721] = c_Body_x[1721];
            n_Body_y[1721] = c_Body_y[1721];
            n_Body_x[1722] = c_Body_x[1722];
            n_Body_y[1722] = c_Body_y[1722];
            n_Body_x[1723] = c_Body_x[1723];
            n_Body_y[1723] = c_Body_y[1723];
            n_Body_x[1724] = c_Body_x[1724];
            n_Body_y[1724] = c_Body_y[1724];
            n_Body_x[1725] = c_Body_x[1725];
            n_Body_y[1725] = c_Body_y[1725];
            n_Body_x[1726] = c_Body_x[1726];
            n_Body_y[1726] = c_Body_y[1726];
            n_Body_x[1727] = c_Body_x[1727];
            n_Body_y[1727] = c_Body_y[1727];
            n_Body_x[1728] = c_Body_x[1728];
            n_Body_y[1728] = c_Body_y[1728];
            n_Body_x[1729] = c_Body_x[1729];
            n_Body_y[1729] = c_Body_y[1729];
            n_Body_x[1730] = c_Body_x[1730];
            n_Body_y[1730] = c_Body_y[1730];
            n_Body_x[1731] = c_Body_x[1731];
            n_Body_y[1731] = c_Body_y[1731];
            n_Body_x[1732] = c_Body_x[1732];
            n_Body_y[1732] = c_Body_y[1732];
            n_Body_x[1733] = c_Body_x[1733];
            n_Body_y[1733] = c_Body_y[1733];
            n_Body_x[1734] = c_Body_x[1734];
            n_Body_y[1734] = c_Body_y[1734];
            n_Body_x[1735] = c_Body_x[1735];
            n_Body_y[1735] = c_Body_y[1735];
            n_Body_x[1736] = c_Body_x[1736];
            n_Body_y[1736] = c_Body_y[1736];
            n_Body_x[1737] = c_Body_x[1737];
            n_Body_y[1737] = c_Body_y[1737];
            n_Body_x[1738] = c_Body_x[1738];
            n_Body_y[1738] = c_Body_y[1738];
            n_Body_x[1739] = c_Body_x[1739];
            n_Body_y[1739] = c_Body_y[1739];
            n_Body_x[1740] = c_Body_x[1740];
            n_Body_y[1740] = c_Body_y[1740];
            n_Body_x[1741] = c_Body_x[1741];
            n_Body_y[1741] = c_Body_y[1741];
            n_Body_x[1742] = c_Body_x[1742];
            n_Body_y[1742] = c_Body_y[1742];
            n_Body_x[1743] = c_Body_x[1743];
            n_Body_y[1743] = c_Body_y[1743];
            n_Body_x[1744] = c_Body_x[1744];
            n_Body_y[1744] = c_Body_y[1744];
            n_Body_x[1745] = c_Body_x[1745];
            n_Body_y[1745] = c_Body_y[1745];
            n_Body_x[1746] = c_Body_x[1746];
            n_Body_y[1746] = c_Body_y[1746];
            n_Body_x[1747] = c_Body_x[1747];
            n_Body_y[1747] = c_Body_y[1747];
            n_Body_x[1748] = c_Body_x[1748];
            n_Body_y[1748] = c_Body_y[1748];
            n_Body_x[1749] = c_Body_x[1749];
            n_Body_y[1749] = c_Body_y[1749];
            n_Body_x[1750] = c_Body_x[1750];
            n_Body_y[1750] = c_Body_y[1750];
            n_Body_x[1751] = c_Body_x[1751];
            n_Body_y[1751] = c_Body_y[1751];
            n_Body_x[1752] = c_Body_x[1752];
            n_Body_y[1752] = c_Body_y[1752];
            n_Body_x[1753] = c_Body_x[1753];
            n_Body_y[1753] = c_Body_y[1753];
            n_Body_x[1754] = c_Body_x[1754];
            n_Body_y[1754] = c_Body_y[1754];
            n_Body_x[1755] = c_Body_x[1755];
            n_Body_y[1755] = c_Body_y[1755];
            n_Body_x[1756] = c_Body_x[1756];
            n_Body_y[1756] = c_Body_y[1756];
            n_Body_x[1757] = c_Body_x[1757];
            n_Body_y[1757] = c_Body_y[1757];
            n_Body_x[1758] = c_Body_x[1758];
            n_Body_y[1758] = c_Body_y[1758];
            n_Body_x[1759] = c_Body_x[1759];
            n_Body_y[1759] = c_Body_y[1759];
            n_Body_x[1760] = c_Body_x[1760];
            n_Body_y[1760] = c_Body_y[1760];
            n_Body_x[1761] = c_Body_x[1761];
            n_Body_y[1761] = c_Body_y[1761];
            n_Body_x[1762] = c_Body_x[1762];
            n_Body_y[1762] = c_Body_y[1762];
            n_Body_x[1763] = c_Body_x[1763];
            n_Body_y[1763] = c_Body_y[1763];
            n_Body_x[1764] = c_Body_x[1764];
            n_Body_y[1764] = c_Body_y[1764];
            n_Body_x[1765] = c_Body_x[1765];
            n_Body_y[1765] = c_Body_y[1765];
            n_Body_x[1766] = c_Body_x[1766];
            n_Body_y[1766] = c_Body_y[1766];
            n_Body_x[1767] = c_Body_x[1767];
            n_Body_y[1767] = c_Body_y[1767];
            n_Body_x[1768] = c_Body_x[1768];
            n_Body_y[1768] = c_Body_y[1768];
            n_Body_x[1769] = c_Body_x[1769];
            n_Body_y[1769] = c_Body_y[1769];
            n_Body_x[1770] = c_Body_x[1770];
            n_Body_y[1770] = c_Body_y[1770];
            n_Body_x[1771] = c_Body_x[1771];
            n_Body_y[1771] = c_Body_y[1771];
            n_Body_x[1772] = c_Body_x[1772];
            n_Body_y[1772] = c_Body_y[1772];
            n_Body_x[1773] = c_Body_x[1773];
            n_Body_y[1773] = c_Body_y[1773];
            n_Body_x[1774] = c_Body_x[1774];
            n_Body_y[1774] = c_Body_y[1774];
            n_Body_x[1775] = c_Body_x[1775];
            n_Body_y[1775] = c_Body_y[1775];
            n_Body_x[1776] = c_Body_x[1776];
            n_Body_y[1776] = c_Body_y[1776];
            n_Body_x[1777] = c_Body_x[1777];
            n_Body_y[1777] = c_Body_y[1777];
            n_Body_x[1778] = c_Body_x[1778];
            n_Body_y[1778] = c_Body_y[1778];
            n_Body_x[1779] = c_Body_x[1779];
            n_Body_y[1779] = c_Body_y[1779];
            n_Body_x[1780] = c_Body_x[1780];
            n_Body_y[1780] = c_Body_y[1780];
            n_Body_x[1781] = c_Body_x[1781];
            n_Body_y[1781] = c_Body_y[1781];
            n_Body_x[1782] = c_Body_x[1782];
            n_Body_y[1782] = c_Body_y[1782];
            n_Body_x[1783] = c_Body_x[1783];
            n_Body_y[1783] = c_Body_y[1783];
            n_Body_x[1784] = c_Body_x[1784];
            n_Body_y[1784] = c_Body_y[1784];
            n_Body_x[1785] = c_Body_x[1785];
            n_Body_y[1785] = c_Body_y[1785];
            n_Body_x[1786] = c_Body_x[1786];
            n_Body_y[1786] = c_Body_y[1786];
            n_Body_x[1787] = c_Body_x[1787];
            n_Body_y[1787] = c_Body_y[1787];
            n_Body_x[1788] = c_Body_x[1788];
            n_Body_y[1788] = c_Body_y[1788];
            n_Body_x[1789] = c_Body_x[1789];
            n_Body_y[1789] = c_Body_y[1789];
            n_Body_x[1790] = c_Body_x[1790];
            n_Body_y[1790] = c_Body_y[1790];
            n_Body_x[1791] = c_Body_x[1791];
            n_Body_y[1791] = c_Body_y[1791];
            n_Body_x[1792] = c_Body_x[1792];
            n_Body_y[1792] = c_Body_y[1792];
            n_Body_x[1793] = c_Body_x[1793];
            n_Body_y[1793] = c_Body_y[1793];
            n_Body_x[1794] = c_Body_x[1794];
            n_Body_y[1794] = c_Body_y[1794];
            n_Body_x[1795] = c_Body_x[1795];
            n_Body_y[1795] = c_Body_y[1795];
            n_Body_x[1796] = c_Body_x[1796];
            n_Body_y[1796] = c_Body_y[1796];
            n_Body_x[1797] = c_Body_x[1797];
            n_Body_y[1797] = c_Body_y[1797];
            n_Body_x[1798] = c_Body_x[1798];
            n_Body_y[1798] = c_Body_y[1798];
            n_Body_x[1799] = c_Body_x[1799];
            n_Body_y[1799] = c_Body_y[1799];
            n_Body_x[1800] = c_Body_x[1800];
            n_Body_y[1800] = c_Body_y[1800];
            n_Body_x[1801] = c_Body_x[1801];
            n_Body_y[1801] = c_Body_y[1801];
            n_Body_x[1802] = c_Body_x[1802];
            n_Body_y[1802] = c_Body_y[1802];
            n_Body_x[1803] = c_Body_x[1803];
            n_Body_y[1803] = c_Body_y[1803];
            n_Body_x[1804] = c_Body_x[1804];
            n_Body_y[1804] = c_Body_y[1804];
            n_Body_x[1805] = c_Body_x[1805];
            n_Body_y[1805] = c_Body_y[1805];
            n_Body_x[1806] = c_Body_x[1806];
            n_Body_y[1806] = c_Body_y[1806];
            n_Body_x[1807] = c_Body_x[1807];
            n_Body_y[1807] = c_Body_y[1807];
            n_Body_x[1808] = c_Body_x[1808];
            n_Body_y[1808] = c_Body_y[1808];
            n_Body_x[1809] = c_Body_x[1809];
            n_Body_y[1809] = c_Body_y[1809];
            n_Body_x[1810] = c_Body_x[1810];
            n_Body_y[1810] = c_Body_y[1810];
            n_Body_x[1811] = c_Body_x[1811];
            n_Body_y[1811] = c_Body_y[1811];
            n_Body_x[1812] = c_Body_x[1812];
            n_Body_y[1812] = c_Body_y[1812];
            n_Body_x[1813] = c_Body_x[1813];
            n_Body_y[1813] = c_Body_y[1813];
            n_Body_x[1814] = c_Body_x[1814];
            n_Body_y[1814] = c_Body_y[1814];
            n_Body_x[1815] = c_Body_x[1815];
            n_Body_y[1815] = c_Body_y[1815];
            n_Body_x[1816] = c_Body_x[1816];
            n_Body_y[1816] = c_Body_y[1816];
            n_Body_x[1817] = c_Body_x[1817];
            n_Body_y[1817] = c_Body_y[1817];
            n_Body_x[1818] = c_Body_x[1818];
            n_Body_y[1818] = c_Body_y[1818];
            n_Body_x[1819] = c_Body_x[1819];
            n_Body_y[1819] = c_Body_y[1819];
            n_Body_x[1820] = c_Body_x[1820];
            n_Body_y[1820] = c_Body_y[1820];
            n_Body_x[1821] = c_Body_x[1821];
            n_Body_y[1821] = c_Body_y[1821];
            n_Body_x[1822] = c_Body_x[1822];
            n_Body_y[1822] = c_Body_y[1822];
            n_Body_x[1823] = c_Body_x[1823];
            n_Body_y[1823] = c_Body_y[1823];
            n_Body_x[1824] = c_Body_x[1824];
            n_Body_y[1824] = c_Body_y[1824];
            n_Body_x[1825] = c_Body_x[1825];
            n_Body_y[1825] = c_Body_y[1825];
            n_Body_x[1826] = c_Body_x[1826];
            n_Body_y[1826] = c_Body_y[1826];
            n_Body_x[1827] = c_Body_x[1827];
            n_Body_y[1827] = c_Body_y[1827];
            n_Body_x[1828] = c_Body_x[1828];
            n_Body_y[1828] = c_Body_y[1828];
            n_Body_x[1829] = c_Body_x[1829];
            n_Body_y[1829] = c_Body_y[1829];
            n_Body_x[1830] = c_Body_x[1830];
            n_Body_y[1830] = c_Body_y[1830];
            n_Body_x[1831] = c_Body_x[1831];
            n_Body_y[1831] = c_Body_y[1831];
            n_Body_x[1832] = c_Body_x[1832];
            n_Body_y[1832] = c_Body_y[1832];
            n_Body_x[1833] = c_Body_x[1833];
            n_Body_y[1833] = c_Body_y[1833];
            n_Body_x[1834] = c_Body_x[1834];
            n_Body_y[1834] = c_Body_y[1834];
            n_Body_x[1835] = c_Body_x[1835];
            n_Body_y[1835] = c_Body_y[1835];
            n_Body_x[1836] = c_Body_x[1836];
            n_Body_y[1836] = c_Body_y[1836];
            n_Body_x[1837] = c_Body_x[1837];
            n_Body_y[1837] = c_Body_y[1837];
            n_Body_x[1838] = c_Body_x[1838];
            n_Body_y[1838] = c_Body_y[1838];
            n_Body_x[1839] = c_Body_x[1839];
            n_Body_y[1839] = c_Body_y[1839];
            n_Body_x[1840] = c_Body_x[1840];
            n_Body_y[1840] = c_Body_y[1840];
            n_Body_x[1841] = c_Body_x[1841];
            n_Body_y[1841] = c_Body_y[1841];
            n_Body_x[1842] = c_Body_x[1842];
            n_Body_y[1842] = c_Body_y[1842];
            n_Body_x[1843] = c_Body_x[1843];
            n_Body_y[1843] = c_Body_y[1843];
            n_Body_x[1844] = c_Body_x[1844];
            n_Body_y[1844] = c_Body_y[1844];
            n_Body_x[1845] = c_Body_x[1845];
            n_Body_y[1845] = c_Body_y[1845];
            n_Body_x[1846] = c_Body_x[1846];
            n_Body_y[1846] = c_Body_y[1846];
            n_Body_x[1847] = c_Body_x[1847];
            n_Body_y[1847] = c_Body_y[1847];
            n_Body_x[1848] = c_Body_x[1848];
            n_Body_y[1848] = c_Body_y[1848];
            n_Body_x[1849] = c_Body_x[1849];
            n_Body_y[1849] = c_Body_y[1849];
            n_Body_x[1850] = c_Body_x[1850];
            n_Body_y[1850] = c_Body_y[1850];
            n_Body_x[1851] = c_Body_x[1851];
            n_Body_y[1851] = c_Body_y[1851];
            n_Body_x[1852] = c_Body_x[1852];
            n_Body_y[1852] = c_Body_y[1852];
            n_Body_x[1853] = c_Body_x[1853];
            n_Body_y[1853] = c_Body_y[1853];
            n_Body_x[1854] = c_Body_x[1854];
            n_Body_y[1854] = c_Body_y[1854];
            n_Body_x[1855] = c_Body_x[1855];
            n_Body_y[1855] = c_Body_y[1855];
            n_Body_x[1856] = c_Body_x[1856];
            n_Body_y[1856] = c_Body_y[1856];
            n_Body_x[1857] = c_Body_x[1857];
            n_Body_y[1857] = c_Body_y[1857];
            n_Body_x[1858] = c_Body_x[1858];
            n_Body_y[1858] = c_Body_y[1858];
            n_Body_x[1859] = c_Body_x[1859];
            n_Body_y[1859] = c_Body_y[1859];
            n_Body_x[1860] = c_Body_x[1860];
            n_Body_y[1860] = c_Body_y[1860];
            n_Body_x[1861] = c_Body_x[1861];
            n_Body_y[1861] = c_Body_y[1861];
            n_Body_x[1862] = c_Body_x[1862];
            n_Body_y[1862] = c_Body_y[1862];
            n_Body_x[1863] = c_Body_x[1863];
            n_Body_y[1863] = c_Body_y[1863];
            n_Body_x[1864] = c_Body_x[1864];
            n_Body_y[1864] = c_Body_y[1864];
            n_Body_x[1865] = c_Body_x[1865];
            n_Body_y[1865] = c_Body_y[1865];
            n_Body_x[1866] = c_Body_x[1866];
            n_Body_y[1866] = c_Body_y[1866];
            n_Body_x[1867] = c_Body_x[1867];
            n_Body_y[1867] = c_Body_y[1867];
            n_Body_x[1868] = c_Body_x[1868];
            n_Body_y[1868] = c_Body_y[1868];
            n_Body_x[1869] = c_Body_x[1869];
            n_Body_y[1869] = c_Body_y[1869];
            n_Body_x[1870] = c_Body_x[1870];
            n_Body_y[1870] = c_Body_y[1870];
            n_Body_x[1871] = c_Body_x[1871];
            n_Body_y[1871] = c_Body_y[1871];
            n_Body_x[1872] = c_Body_x[1872];
            n_Body_y[1872] = c_Body_y[1872];
            n_Body_x[1873] = c_Body_x[1873];
            n_Body_y[1873] = c_Body_y[1873];
            n_Body_x[1874] = c_Body_x[1874];
            n_Body_y[1874] = c_Body_y[1874];
            n_Body_x[1875] = c_Body_x[1875];
            n_Body_y[1875] = c_Body_y[1875];
            n_Body_x[1876] = c_Body_x[1876];
            n_Body_y[1876] = c_Body_y[1876];
            n_Body_x[1877] = c_Body_x[1877];
            n_Body_y[1877] = c_Body_y[1877];
            n_Body_x[1878] = c_Body_x[1878];
            n_Body_y[1878] = c_Body_y[1878];
            n_Body_x[1879] = c_Body_x[1879];
            n_Body_y[1879] = c_Body_y[1879];
            n_Body_x[1880] = c_Body_x[1880];
            n_Body_y[1880] = c_Body_y[1880];
            n_Body_x[1881] = c_Body_x[1881];
            n_Body_y[1881] = c_Body_y[1881];
            n_Body_x[1882] = c_Body_x[1882];
            n_Body_y[1882] = c_Body_y[1882];
            n_Body_x[1883] = c_Body_x[1883];
            n_Body_y[1883] = c_Body_y[1883];
            n_Body_x[1884] = c_Body_x[1884];
            n_Body_y[1884] = c_Body_y[1884];
            n_Body_x[1885] = c_Body_x[1885];
            n_Body_y[1885] = c_Body_y[1885];
            n_Body_x[1886] = c_Body_x[1886];
            n_Body_y[1886] = c_Body_y[1886];
            n_Body_x[1887] = c_Body_x[1887];
            n_Body_y[1887] = c_Body_y[1887];
            n_Body_x[1888] = c_Body_x[1888];
            n_Body_y[1888] = c_Body_y[1888];
            n_Body_x[1889] = c_Body_x[1889];
            n_Body_y[1889] = c_Body_y[1889];
            n_Body_x[1890] = c_Body_x[1890];
            n_Body_y[1890] = c_Body_y[1890];
            n_Body_x[1891] = c_Body_x[1891];
            n_Body_y[1891] = c_Body_y[1891];
            n_Body_x[1892] = c_Body_x[1892];
            n_Body_y[1892] = c_Body_y[1892];
            n_Body_x[1893] = c_Body_x[1893];
            n_Body_y[1893] = c_Body_y[1893];
            n_Body_x[1894] = c_Body_x[1894];
            n_Body_y[1894] = c_Body_y[1894];
            n_Body_x[1895] = c_Body_x[1895];
            n_Body_y[1895] = c_Body_y[1895];
            n_Body_x[1896] = c_Body_x[1896];
            n_Body_y[1896] = c_Body_y[1896];
            n_Body_x[1897] = c_Body_x[1897];
            n_Body_y[1897] = c_Body_y[1897];
            n_Body_x[1898] = c_Body_x[1898];
            n_Body_y[1898] = c_Body_y[1898];
            n_Body_x[1899] = c_Body_x[1899];
            n_Body_y[1899] = c_Body_y[1899];
            n_Body_x[1900] = c_Body_x[1900];
            n_Body_y[1900] = c_Body_y[1900];
            n_Body_x[1901] = c_Body_x[1901];
            n_Body_y[1901] = c_Body_y[1901];
            n_Body_x[1902] = c_Body_x[1902];
            n_Body_y[1902] = c_Body_y[1902];
            n_Body_x[1903] = c_Body_x[1903];
            n_Body_y[1903] = c_Body_y[1903];
            n_Body_x[1904] = c_Body_x[1904];
            n_Body_y[1904] = c_Body_y[1904];
            n_Body_x[1905] = c_Body_x[1905];
            n_Body_y[1905] = c_Body_y[1905];
            n_Body_x[1906] = c_Body_x[1906];
            n_Body_y[1906] = c_Body_y[1906];
            n_Body_x[1907] = c_Body_x[1907];
            n_Body_y[1907] = c_Body_y[1907];
            n_Body_x[1908] = c_Body_x[1908];
            n_Body_y[1908] = c_Body_y[1908];
            n_Body_x[1909] = c_Body_x[1909];
            n_Body_y[1909] = c_Body_y[1909];
            n_Body_x[1910] = c_Body_x[1910];
            n_Body_y[1910] = c_Body_y[1910];
            n_Body_x[1911] = c_Body_x[1911];
            n_Body_y[1911] = c_Body_y[1911];
            n_Body_x[1912] = c_Body_x[1912];
            n_Body_y[1912] = c_Body_y[1912];
            n_Body_x[1913] = c_Body_x[1913];
            n_Body_y[1913] = c_Body_y[1913];
            n_Body_x[1914] = c_Body_x[1914];
            n_Body_y[1914] = c_Body_y[1914];
            n_Body_x[1915] = c_Body_x[1915];
            n_Body_y[1915] = c_Body_y[1915];
            n_Body_x[1916] = c_Body_x[1916];
            n_Body_y[1916] = c_Body_y[1916];
            n_Body_x[1917] = c_Body_x[1917];
            n_Body_y[1917] = c_Body_y[1917];
            n_Body_x[1918] = c_Body_x[1918];
            n_Body_y[1918] = c_Body_y[1918];
            n_Body_x[1919] = c_Body_x[1919];
            n_Body_y[1919] = c_Body_y[1919];
            n_Body_x[1920] = c_Body_x[1920];
            n_Body_y[1920] = c_Body_y[1920];
            n_Body_x[1921] = c_Body_x[1921];
            n_Body_y[1921] = c_Body_y[1921];
            n_Body_x[1922] = c_Body_x[1922];
            n_Body_y[1922] = c_Body_y[1922];
            n_Body_x[1923] = c_Body_x[1923];
            n_Body_y[1923] = c_Body_y[1923];
            n_Body_x[1924] = c_Body_x[1924];
            n_Body_y[1924] = c_Body_y[1924];
            n_Body_x[1925] = c_Body_x[1925];
            n_Body_y[1925] = c_Body_y[1925];
            n_Body_x[1926] = c_Body_x[1926];
            n_Body_y[1926] = c_Body_y[1926];
            n_Body_x[1927] = c_Body_x[1927];
            n_Body_y[1927] = c_Body_y[1927];
            n_Body_x[1928] = c_Body_x[1928];
            n_Body_y[1928] = c_Body_y[1928];
            n_Body_x[1929] = c_Body_x[1929];
            n_Body_y[1929] = c_Body_y[1929];
            n_Body_x[1930] = c_Body_x[1930];
            n_Body_y[1930] = c_Body_y[1930];
            n_Body_x[1931] = c_Body_x[1931];
            n_Body_y[1931] = c_Body_y[1931];
            n_Body_x[1932] = c_Body_x[1932];
            n_Body_y[1932] = c_Body_y[1932];
            n_Body_x[1933] = c_Body_x[1933];
            n_Body_y[1933] = c_Body_y[1933];
            n_Body_x[1934] = c_Body_x[1934];
            n_Body_y[1934] = c_Body_y[1934];
            n_Body_x[1935] = c_Body_x[1935];
            n_Body_y[1935] = c_Body_y[1935];
            n_Body_x[1936] = c_Body_x[1936];
            n_Body_y[1936] = c_Body_y[1936];
            n_Body_x[1937] = c_Body_x[1937];
            n_Body_y[1937] = c_Body_y[1937];
            n_Body_x[1938] = c_Body_x[1938];
            n_Body_y[1938] = c_Body_y[1938];
            n_Body_x[1939] = c_Body_x[1939];
            n_Body_y[1939] = c_Body_y[1939];
            n_Body_x[1940] = c_Body_x[1940];
            n_Body_y[1940] = c_Body_y[1940];
            n_Body_x[1941] = c_Body_x[1941];
            n_Body_y[1941] = c_Body_y[1941];
            n_Body_x[1942] = c_Body_x[1942];
            n_Body_y[1942] = c_Body_y[1942];
            n_Body_x[1943] = c_Body_x[1943];
            n_Body_y[1943] = c_Body_y[1943];
            n_Body_x[1944] = c_Body_x[1944];
            n_Body_y[1944] = c_Body_y[1944];
            n_Body_x[1945] = c_Body_x[1945];
            n_Body_y[1945] = c_Body_y[1945];
            n_Body_x[1946] = c_Body_x[1946];
            n_Body_y[1946] = c_Body_y[1946];
            n_Body_x[1947] = c_Body_x[1947];
            n_Body_y[1947] = c_Body_y[1947];
            n_Body_x[1948] = c_Body_x[1948];
            n_Body_y[1948] = c_Body_y[1948];
            n_Body_x[1949] = c_Body_x[1949];
            n_Body_y[1949] = c_Body_y[1949];
            n_Body_x[1950] = c_Body_x[1950];
            n_Body_y[1950] = c_Body_y[1950];
            n_Body_x[1951] = c_Body_x[1951];
            n_Body_y[1951] = c_Body_y[1951];
            n_Body_x[1952] = c_Body_x[1952];
            n_Body_y[1952] = c_Body_y[1952];
            n_Body_x[1953] = c_Body_x[1953];
            n_Body_y[1953] = c_Body_y[1953];
            n_Body_x[1954] = c_Body_x[1954];
            n_Body_y[1954] = c_Body_y[1954];
            n_Body_x[1955] = c_Body_x[1955];
            n_Body_y[1955] = c_Body_y[1955];
            n_Body_x[1956] = c_Body_x[1956];
            n_Body_y[1956] = c_Body_y[1956];
            n_Body_x[1957] = c_Body_x[1957];
            n_Body_y[1957] = c_Body_y[1957];
            n_Body_x[1958] = c_Body_x[1958];
            n_Body_y[1958] = c_Body_y[1958];
            n_Body_x[1959] = c_Body_x[1959];
            n_Body_y[1959] = c_Body_y[1959];
            n_Body_x[1960] = c_Body_x[1960];
            n_Body_y[1960] = c_Body_y[1960];
            n_Body_x[1961] = c_Body_x[1961];
            n_Body_y[1961] = c_Body_y[1961];
            n_Body_x[1962] = c_Body_x[1962];
            n_Body_y[1962] = c_Body_y[1962];
            n_Body_x[1963] = c_Body_x[1963];
            n_Body_y[1963] = c_Body_y[1963];
            n_Body_x[1964] = c_Body_x[1964];
            n_Body_y[1964] = c_Body_y[1964];
            n_Body_x[1965] = c_Body_x[1965];
            n_Body_y[1965] = c_Body_y[1965];
            n_Body_x[1966] = c_Body_x[1966];
            n_Body_y[1966] = c_Body_y[1966];
            n_Body_x[1967] = c_Body_x[1967];
            n_Body_y[1967] = c_Body_y[1967];
            n_Body_x[1968] = c_Body_x[1968];
            n_Body_y[1968] = c_Body_y[1968];
            n_Body_x[1969] = c_Body_x[1969];
            n_Body_y[1969] = c_Body_y[1969];
            n_Body_x[1970] = c_Body_x[1970];
            n_Body_y[1970] = c_Body_y[1970];
            n_Body_x[1971] = c_Body_x[1971];
            n_Body_y[1971] = c_Body_y[1971];
            n_Body_x[1972] = c_Body_x[1972];
            n_Body_y[1972] = c_Body_y[1972];
            n_Body_x[1973] = c_Body_x[1973];
            n_Body_y[1973] = c_Body_y[1973];
            n_Body_x[1974] = c_Body_x[1974];
            n_Body_y[1974] = c_Body_y[1974];
            n_Body_x[1975] = c_Body_x[1975];
            n_Body_y[1975] = c_Body_y[1975];
            n_Body_x[1976] = c_Body_x[1976];
            n_Body_y[1976] = c_Body_y[1976];
            n_Body_x[1977] = c_Body_x[1977];
            n_Body_y[1977] = c_Body_y[1977];
            n_Body_x[1978] = c_Body_x[1978];
            n_Body_y[1978] = c_Body_y[1978];
            n_Body_x[1979] = c_Body_x[1979];
            n_Body_y[1979] = c_Body_y[1979];
            n_Body_x[1980] = c_Body_x[1980];
            n_Body_y[1980] = c_Body_y[1980];
            n_Body_x[1981] = c_Body_x[1981];
            n_Body_y[1981] = c_Body_y[1981];
            n_Body_x[1982] = c_Body_x[1982];
            n_Body_y[1982] = c_Body_y[1982];
            n_Body_x[1983] = c_Body_x[1983];
            n_Body_y[1983] = c_Body_y[1983];
            n_Body_x[1984] = c_Body_x[1984];
            n_Body_y[1984] = c_Body_y[1984];
            n_Body_x[1985] = c_Body_x[1985];
            n_Body_y[1985] = c_Body_y[1985];
            n_Body_x[1986] = c_Body_x[1986];
            n_Body_y[1986] = c_Body_y[1986];
            n_Body_x[1987] = c_Body_x[1987];
            n_Body_y[1987] = c_Body_y[1987];
            n_Body_x[1988] = c_Body_x[1988];
            n_Body_y[1988] = c_Body_y[1988];
            n_Body_x[1989] = c_Body_x[1989];
            n_Body_y[1989] = c_Body_y[1989];
            n_Body_x[1990] = c_Body_x[1990];
            n_Body_y[1990] = c_Body_y[1990];
            n_Body_x[1991] = c_Body_x[1991];
            n_Body_y[1991] = c_Body_y[1991];
            n_Body_x[1992] = c_Body_x[1992];
            n_Body_y[1992] = c_Body_y[1992];
            n_Body_x[1993] = c_Body_x[1993];
            n_Body_y[1993] = c_Body_y[1993];
            n_Body_x[1994] = c_Body_x[1994];
            n_Body_y[1994] = c_Body_y[1994];
            n_Body_x[1995] = c_Body_x[1995];
            n_Body_y[1995] = c_Body_y[1995];
            n_Body_x[1996] = c_Body_x[1996];
            n_Body_y[1996] = c_Body_y[1996];
            n_Body_x[1997] = c_Body_x[1997];
            n_Body_y[1997] = c_Body_y[1997];
            n_Body_x[1998] = c_Body_x[1998];
            n_Body_y[1998] = c_Body_y[1998];
            n_Body_x[1999] = c_Body_x[1999];
            n_Body_y[1999] = c_Body_y[1999];
            n_Body_x[2000] = c_Body_x[2000];
            n_Body_y[2000] = c_Body_y[2000];
            n_Body_x[2001] = c_Body_x[2001];
            n_Body_y[2001] = c_Body_y[2001];
            n_Body_x[2002] = c_Body_x[2002];
            n_Body_y[2002] = c_Body_y[2002];
            n_Body_x[2003] = c_Body_x[2003];
            n_Body_y[2003] = c_Body_y[2003];
            n_Body_x[2004] = c_Body_x[2004];
            n_Body_y[2004] = c_Body_y[2004];
            n_Body_x[2005] = c_Body_x[2005];
            n_Body_y[2005] = c_Body_y[2005];
            n_Body_x[2006] = c_Body_x[2006];
            n_Body_y[2006] = c_Body_y[2006];
            n_Body_x[2007] = c_Body_x[2007];
            n_Body_y[2007] = c_Body_y[2007];
            n_Body_x[2008] = c_Body_x[2008];
            n_Body_y[2008] = c_Body_y[2008];
            n_Body_x[2009] = c_Body_x[2009];
            n_Body_y[2009] = c_Body_y[2009];
            n_Body_x[2010] = c_Body_x[2010];
            n_Body_y[2010] = c_Body_y[2010];
            n_Body_x[2011] = c_Body_x[2011];
            n_Body_y[2011] = c_Body_y[2011];
            n_Body_x[2012] = c_Body_x[2012];
            n_Body_y[2012] = c_Body_y[2012];
            n_Body_x[2013] = c_Body_x[2013];
            n_Body_y[2013] = c_Body_y[2013];
            n_Body_x[2014] = c_Body_x[2014];
            n_Body_y[2014] = c_Body_y[2014];
            n_Body_x[2015] = c_Body_x[2015];
            n_Body_y[2015] = c_Body_y[2015];
            n_Body_x[2016] = c_Body_x[2016];
            n_Body_y[2016] = c_Body_y[2016];
            n_Body_x[2017] = c_Body_x[2017];
            n_Body_y[2017] = c_Body_y[2017];
            n_Body_x[2018] = c_Body_x[2018];
            n_Body_y[2018] = c_Body_y[2018];
            n_Body_x[2019] = c_Body_x[2019];
            n_Body_y[2019] = c_Body_y[2019];
            n_Body_x[2020] = c_Body_x[2020];
            n_Body_y[2020] = c_Body_y[2020];
            n_Body_x[2021] = c_Body_x[2021];
            n_Body_y[2021] = c_Body_y[2021];
            n_Body_x[2022] = c_Body_x[2022];
            n_Body_y[2022] = c_Body_y[2022];
            n_Body_x[2023] = c_Body_x[2023];
            n_Body_y[2023] = c_Body_y[2023];
            n_Body_x[2024] = c_Body_x[2024];
            n_Body_y[2024] = c_Body_y[2024];
            n_Body_x[2025] = c_Body_x[2025];
            n_Body_y[2025] = c_Body_y[2025];
            n_Body_x[2026] = c_Body_x[2026];
            n_Body_y[2026] = c_Body_y[2026];
            n_Body_x[2027] = c_Body_x[2027];
            n_Body_y[2027] = c_Body_y[2027];
            n_Body_x[2028] = c_Body_x[2028];
            n_Body_y[2028] = c_Body_y[2028];
            n_Body_x[2029] = c_Body_x[2029];
            n_Body_y[2029] = c_Body_y[2029];
            n_Body_x[2030] = c_Body_x[2030];
            n_Body_y[2030] = c_Body_y[2030];
            n_Body_x[2031] = c_Body_x[2031];
            n_Body_y[2031] = c_Body_y[2031];
            n_Body_x[2032] = c_Body_x[2032];
            n_Body_y[2032] = c_Body_y[2032];
            n_Body_x[2033] = c_Body_x[2033];
            n_Body_y[2033] = c_Body_y[2033];
            n_Body_x[2034] = c_Body_x[2034];
            n_Body_y[2034] = c_Body_y[2034];
            n_Body_x[2035] = c_Body_x[2035];
            n_Body_y[2035] = c_Body_y[2035];
            n_Body_x[2036] = c_Body_x[2036];
            n_Body_y[2036] = c_Body_y[2036];
            n_Body_x[2037] = c_Body_x[2037];
            n_Body_y[2037] = c_Body_y[2037];
            n_Body_x[2038] = c_Body_x[2038];
            n_Body_y[2038] = c_Body_y[2038];
            n_Body_x[2039] = c_Body_x[2039];
            n_Body_y[2039] = c_Body_y[2039];
            n_Body_x[2040] = c_Body_x[2040];
            n_Body_y[2040] = c_Body_y[2040];
            n_Body_x[2041] = c_Body_x[2041];
            n_Body_y[2041] = c_Body_y[2041];
            n_Body_x[2042] = c_Body_x[2042];
            n_Body_y[2042] = c_Body_y[2042];
            n_Body_x[2043] = c_Body_x[2043];
            n_Body_y[2043] = c_Body_y[2043];
            n_Body_x[2044] = c_Body_x[2044];
            n_Body_y[2044] = c_Body_y[2044];
            n_Body_x[2045] = c_Body_x[2045];
            n_Body_y[2045] = c_Body_y[2045];
            n_Body_x[2046] = c_Body_x[2046];
            n_Body_y[2046] = c_Body_y[2046];
            n_Body_x[2047] = c_Body_x[2047];
            n_Body_y[2047] = c_Body_y[2047];
            n_Body_x[2048] = c_Body_x[2048];
            n_Body_y[2048] = c_Body_y[2048];
            n_Body_x[2049] = c_Body_x[2049];
            n_Body_y[2049] = c_Body_y[2049];
            n_Body_x[2050] = c_Body_x[2050];
            n_Body_y[2050] = c_Body_y[2050];
            n_Body_x[2051] = c_Body_x[2051];
            n_Body_y[2051] = c_Body_y[2051];
            n_Body_x[2052] = c_Body_x[2052];
            n_Body_y[2052] = c_Body_y[2052];
            n_Body_x[2053] = c_Body_x[2053];
            n_Body_y[2053] = c_Body_y[2053];
            n_Body_x[2054] = c_Body_x[2054];
            n_Body_y[2054] = c_Body_y[2054];
            n_Body_x[2055] = c_Body_x[2055];
            n_Body_y[2055] = c_Body_y[2055];
            n_Body_x[2056] = c_Body_x[2056];
            n_Body_y[2056] = c_Body_y[2056];
            n_Body_x[2057] = c_Body_x[2057];
            n_Body_y[2057] = c_Body_y[2057];
            n_Body_x[2058] = c_Body_x[2058];
            n_Body_y[2058] = c_Body_y[2058];
            n_Body_x[2059] = c_Body_x[2059];
            n_Body_y[2059] = c_Body_y[2059];
            n_Body_x[2060] = c_Body_x[2060];
            n_Body_y[2060] = c_Body_y[2060];
            n_Body_x[2061] = c_Body_x[2061];
            n_Body_y[2061] = c_Body_y[2061];
            n_Body_x[2062] = c_Body_x[2062];
            n_Body_y[2062] = c_Body_y[2062];
            n_Body_x[2063] = c_Body_x[2063];
            n_Body_y[2063] = c_Body_y[2063];
            n_Body_x[2064] = c_Body_x[2064];
            n_Body_y[2064] = c_Body_y[2064];
            n_Body_x[2065] = c_Body_x[2065];
            n_Body_y[2065] = c_Body_y[2065];
            n_Body_x[2066] = c_Body_x[2066];
            n_Body_y[2066] = c_Body_y[2066];
            n_Body_x[2067] = c_Body_x[2067];
            n_Body_y[2067] = c_Body_y[2067];
            n_Body_x[2068] = c_Body_x[2068];
            n_Body_y[2068] = c_Body_y[2068];
            n_Body_x[2069] = c_Body_x[2069];
            n_Body_y[2069] = c_Body_y[2069];
            n_Body_x[2070] = c_Body_x[2070];
            n_Body_y[2070] = c_Body_y[2070];
            n_Body_x[2071] = c_Body_x[2071];
            n_Body_y[2071] = c_Body_y[2071];
            n_Body_x[2072] = c_Body_x[2072];
            n_Body_y[2072] = c_Body_y[2072];
            n_Body_x[2073] = c_Body_x[2073];
            n_Body_y[2073] = c_Body_y[2073];
            n_Body_x[2074] = c_Body_x[2074];
            n_Body_y[2074] = c_Body_y[2074];
            n_Body_x[2075] = c_Body_x[2075];
            n_Body_y[2075] = c_Body_y[2075];
            n_Body_x[2076] = c_Body_x[2076];
            n_Body_y[2076] = c_Body_y[2076];
            n_Body_x[2077] = c_Body_x[2077];
            n_Body_y[2077] = c_Body_y[2077];
            n_Body_x[2078] = c_Body_x[2078];
            n_Body_y[2078] = c_Body_y[2078];
            n_Body_x[2079] = c_Body_x[2079];
            n_Body_y[2079] = c_Body_y[2079];
            n_Body_x[2080] = c_Body_x[2080];
            n_Body_y[2080] = c_Body_y[2080];
            n_Body_x[2081] = c_Body_x[2081];
            n_Body_y[2081] = c_Body_y[2081];
            n_Body_x[2082] = c_Body_x[2082];
            n_Body_y[2082] = c_Body_y[2082];
            n_Body_x[2083] = c_Body_x[2083];
            n_Body_y[2083] = c_Body_y[2083];
            n_Body_x[2084] = c_Body_x[2084];
            n_Body_y[2084] = c_Body_y[2084];
            n_Body_x[2085] = c_Body_x[2085];
            n_Body_y[2085] = c_Body_y[2085];
            n_Body_x[2086] = c_Body_x[2086];
            n_Body_y[2086] = c_Body_y[2086];
            n_Body_x[2087] = c_Body_x[2087];
            n_Body_y[2087] = c_Body_y[2087];
            n_Body_x[2088] = c_Body_x[2088];
            n_Body_y[2088] = c_Body_y[2088];
            n_Body_x[2089] = c_Body_x[2089];
            n_Body_y[2089] = c_Body_y[2089];
            n_Body_x[2090] = c_Body_x[2090];
            n_Body_y[2090] = c_Body_y[2090];
            n_Body_x[2091] = c_Body_x[2091];
            n_Body_y[2091] = c_Body_y[2091];
            n_Body_x[2092] = c_Body_x[2092];
            n_Body_y[2092] = c_Body_y[2092];
            n_Body_x[2093] = c_Body_x[2093];
            n_Body_y[2093] = c_Body_y[2093];
            n_Body_x[2094] = c_Body_x[2094];
            n_Body_y[2094] = c_Body_y[2094];
            n_Body_x[2095] = c_Body_x[2095];
            n_Body_y[2095] = c_Body_y[2095];
            n_Body_x[2096] = c_Body_x[2096];
            n_Body_y[2096] = c_Body_y[2096];
            n_Body_x[2097] = c_Body_x[2097];
            n_Body_y[2097] = c_Body_y[2097];
            n_Body_x[2098] = c_Body_x[2098];
            n_Body_y[2098] = c_Body_y[2098];
            n_Body_x[2099] = c_Body_x[2099];
            n_Body_y[2099] = c_Body_y[2099];
            n_Body_x[2100] = c_Body_x[2100];
            n_Body_y[2100] = c_Body_y[2100];
            n_Body_x[2101] = c_Body_x[2101];
            n_Body_y[2101] = c_Body_y[2101];
            n_Body_x[2102] = c_Body_x[2102];
            n_Body_y[2102] = c_Body_y[2102];
            n_Body_x[2103] = c_Body_x[2103];
            n_Body_y[2103] = c_Body_y[2103];
            n_Body_x[2104] = c_Body_x[2104];
            n_Body_y[2104] = c_Body_y[2104];
            n_Body_x[2105] = c_Body_x[2105];
            n_Body_y[2105] = c_Body_y[2105];
            n_Body_x[2106] = c_Body_x[2106];
            n_Body_y[2106] = c_Body_y[2106];
            n_Body_x[2107] = c_Body_x[2107];
            n_Body_y[2107] = c_Body_y[2107];
            n_Body_x[2108] = c_Body_x[2108];
            n_Body_y[2108] = c_Body_y[2108];
            n_Body_x[2109] = c_Body_x[2109];
            n_Body_y[2109] = c_Body_y[2109];
            n_Body_x[2110] = c_Body_x[2110];
            n_Body_y[2110] = c_Body_y[2110];
            n_Body_x[2111] = c_Body_x[2111];
            n_Body_y[2111] = c_Body_y[2111];
            n_Body_x[2112] = c_Body_x[2112];
            n_Body_y[2112] = c_Body_y[2112];
            n_Body_x[2113] = c_Body_x[2113];
            n_Body_y[2113] = c_Body_y[2113];
            n_Body_x[2114] = c_Body_x[2114];
            n_Body_y[2114] = c_Body_y[2114];
            n_Body_x[2115] = c_Body_x[2115];
            n_Body_y[2115] = c_Body_y[2115];
            n_Body_x[2116] = c_Body_x[2116];
            n_Body_y[2116] = c_Body_y[2116];
            n_Body_x[2117] = c_Body_x[2117];
            n_Body_y[2117] = c_Body_y[2117];
            n_Body_x[2118] = c_Body_x[2118];
            n_Body_y[2118] = c_Body_y[2118];
            n_Body_x[2119] = c_Body_x[2119];
            n_Body_y[2119] = c_Body_y[2119];
            n_Body_x[2120] = c_Body_x[2120];
            n_Body_y[2120] = c_Body_y[2120];
            n_Body_x[2121] = c_Body_x[2121];
            n_Body_y[2121] = c_Body_y[2121];
            n_Body_x[2122] = c_Body_x[2122];
            n_Body_y[2122] = c_Body_y[2122];
            n_Body_x[2123] = c_Body_x[2123];
            n_Body_y[2123] = c_Body_y[2123];
            n_Body_x[2124] = c_Body_x[2124];
            n_Body_y[2124] = c_Body_y[2124];
            n_Body_x[2125] = c_Body_x[2125];
            n_Body_y[2125] = c_Body_y[2125];
            n_Body_x[2126] = c_Body_x[2126];
            n_Body_y[2126] = c_Body_y[2126];
            n_Body_x[2127] = c_Body_x[2127];
            n_Body_y[2127] = c_Body_y[2127];
            n_Body_x[2128] = c_Body_x[2128];
            n_Body_y[2128] = c_Body_y[2128];
            n_Body_x[2129] = c_Body_x[2129];
            n_Body_y[2129] = c_Body_y[2129];
            n_Body_x[2130] = c_Body_x[2130];
            n_Body_y[2130] = c_Body_y[2130];
            n_Body_x[2131] = c_Body_x[2131];
            n_Body_y[2131] = c_Body_y[2131];
            n_Body_x[2132] = c_Body_x[2132];
            n_Body_y[2132] = c_Body_y[2132];
            n_Body_x[2133] = c_Body_x[2133];
            n_Body_y[2133] = c_Body_y[2133];
            n_Body_x[2134] = c_Body_x[2134];
            n_Body_y[2134] = c_Body_y[2134];
            n_Body_x[2135] = c_Body_x[2135];
            n_Body_y[2135] = c_Body_y[2135];
            n_Body_x[2136] = c_Body_x[2136];
            n_Body_y[2136] = c_Body_y[2136];
            n_Body_x[2137] = c_Body_x[2137];
            n_Body_y[2137] = c_Body_y[2137];
            n_Body_x[2138] = c_Body_x[2138];
            n_Body_y[2138] = c_Body_y[2138];
            n_Body_x[2139] = c_Body_x[2139];
            n_Body_y[2139] = c_Body_y[2139];
            n_Body_x[2140] = c_Body_x[2140];
            n_Body_y[2140] = c_Body_y[2140];
            n_Body_x[2141] = c_Body_x[2141];
            n_Body_y[2141] = c_Body_y[2141];
            n_Body_x[2142] = c_Body_x[2142];
            n_Body_y[2142] = c_Body_y[2142];
            n_Body_x[2143] = c_Body_x[2143];
            n_Body_y[2143] = c_Body_y[2143];
            n_Body_x[2144] = c_Body_x[2144];
            n_Body_y[2144] = c_Body_y[2144];
            n_Body_x[2145] = c_Body_x[2145];
            n_Body_y[2145] = c_Body_y[2145];
            n_Body_x[2146] = c_Body_x[2146];
            n_Body_y[2146] = c_Body_y[2146];
            n_Body_x[2147] = c_Body_x[2147];
            n_Body_y[2147] = c_Body_y[2147];
            n_Body_x[2148] = c_Body_x[2148];
            n_Body_y[2148] = c_Body_y[2148];
            n_Body_x[2149] = c_Body_x[2149];
            n_Body_y[2149] = c_Body_y[2149];
            n_Body_x[2150] = c_Body_x[2150];
            n_Body_y[2150] = c_Body_y[2150];
            n_Body_x[2151] = c_Body_x[2151];
            n_Body_y[2151] = c_Body_y[2151];
            n_Body_x[2152] = c_Body_x[2152];
            n_Body_y[2152] = c_Body_y[2152];
            n_Body_x[2153] = c_Body_x[2153];
            n_Body_y[2153] = c_Body_y[2153];
            n_Body_x[2154] = c_Body_x[2154];
            n_Body_y[2154] = c_Body_y[2154];
            n_Body_x[2155] = c_Body_x[2155];
            n_Body_y[2155] = c_Body_y[2155];
            n_Body_x[2156] = c_Body_x[2156];
            n_Body_y[2156] = c_Body_y[2156];
            n_Body_x[2157] = c_Body_x[2157];
            n_Body_y[2157] = c_Body_y[2157];
            n_Body_x[2158] = c_Body_x[2158];
            n_Body_y[2158] = c_Body_y[2158];
            n_Body_x[2159] = c_Body_x[2159];
            n_Body_y[2159] = c_Body_y[2159];
            n_Body_x[2160] = c_Body_x[2160];
            n_Body_y[2160] = c_Body_y[2160];
            n_Body_x[2161] = c_Body_x[2161];
            n_Body_y[2161] = c_Body_y[2161];
            n_Body_x[2162] = c_Body_x[2162];
            n_Body_y[2162] = c_Body_y[2162];
            n_Body_x[2163] = c_Body_x[2163];
            n_Body_y[2163] = c_Body_y[2163];
            n_Body_x[2164] = c_Body_x[2164];
            n_Body_y[2164] = c_Body_y[2164];
            n_Body_x[2165] = c_Body_x[2165];
            n_Body_y[2165] = c_Body_y[2165];
            n_Body_x[2166] = c_Body_x[2166];
            n_Body_y[2166] = c_Body_y[2166];
            n_Body_x[2167] = c_Body_x[2167];
            n_Body_y[2167] = c_Body_y[2167];
            n_Body_x[2168] = c_Body_x[2168];
            n_Body_y[2168] = c_Body_y[2168];
            n_Body_x[2169] = c_Body_x[2169];
            n_Body_y[2169] = c_Body_y[2169];
            n_Body_x[2170] = c_Body_x[2170];
            n_Body_y[2170] = c_Body_y[2170];
            n_Body_x[2171] = c_Body_x[2171];
            n_Body_y[2171] = c_Body_y[2171];
            n_Body_x[2172] = c_Body_x[2172];
            n_Body_y[2172] = c_Body_y[2172];
            n_Body_x[2173] = c_Body_x[2173];
            n_Body_y[2173] = c_Body_y[2173];
            n_Body_x[2174] = c_Body_x[2174];
            n_Body_y[2174] = c_Body_y[2174];
            n_Body_x[2175] = c_Body_x[2175];
            n_Body_y[2175] = c_Body_y[2175];
            n_Body_x[2176] = c_Body_x[2176];
            n_Body_y[2176] = c_Body_y[2176];
            n_Body_x[2177] = c_Body_x[2177];
            n_Body_y[2177] = c_Body_y[2177];
            n_Body_x[2178] = c_Body_x[2178];
            n_Body_y[2178] = c_Body_y[2178];
            n_Body_x[2179] = c_Body_x[2179];
            n_Body_y[2179] = c_Body_y[2179];
            n_Body_x[2180] = c_Body_x[2180];
            n_Body_y[2180] = c_Body_y[2180];
            n_Body_x[2181] = c_Body_x[2181];
            n_Body_y[2181] = c_Body_y[2181];
            n_Body_x[2182] = c_Body_x[2182];
            n_Body_y[2182] = c_Body_y[2182];
            n_Body_x[2183] = c_Body_x[2183];
            n_Body_y[2183] = c_Body_y[2183];
            n_Body_x[2184] = c_Body_x[2184];
            n_Body_y[2184] = c_Body_y[2184];
            n_Body_x[2185] = c_Body_x[2185];
            n_Body_y[2185] = c_Body_y[2185];
            n_Body_x[2186] = c_Body_x[2186];
            n_Body_y[2186] = c_Body_y[2186];
            n_Body_x[2187] = c_Body_x[2187];
            n_Body_y[2187] = c_Body_y[2187];
            n_Body_x[2188] = c_Body_x[2188];
            n_Body_y[2188] = c_Body_y[2188];
            n_Body_x[2189] = c_Body_x[2189];
            n_Body_y[2189] = c_Body_y[2189];
            n_Body_x[2190] = c_Body_x[2190];
            n_Body_y[2190] = c_Body_y[2190];
            n_Body_x[2191] = c_Body_x[2191];
            n_Body_y[2191] = c_Body_y[2191];
            n_Body_x[2192] = c_Body_x[2192];
            n_Body_y[2192] = c_Body_y[2192];
            n_Body_x[2193] = c_Body_x[2193];
            n_Body_y[2193] = c_Body_y[2193];
            n_Body_x[2194] = c_Body_x[2194];
            n_Body_y[2194] = c_Body_y[2194];
            n_Body_x[2195] = c_Body_x[2195];
            n_Body_y[2195] = c_Body_y[2195];
            n_Body_x[2196] = c_Body_x[2196];
            n_Body_y[2196] = c_Body_y[2196];
            n_Body_x[2197] = c_Body_x[2197];
            n_Body_y[2197] = c_Body_y[2197];
            n_Body_x[2198] = c_Body_x[2198];
            n_Body_y[2198] = c_Body_y[2198];
            n_Body_x[2199] = c_Body_x[2199];
            n_Body_y[2199] = c_Body_y[2199];
            n_Body_x[2200] = c_Body_x[2200];
            n_Body_y[2200] = c_Body_y[2200];
            n_Body_x[2201] = c_Body_x[2201];
            n_Body_y[2201] = c_Body_y[2201];
            n_Body_x[2202] = c_Body_x[2202];
            n_Body_y[2202] = c_Body_y[2202];
            n_Body_x[2203] = c_Body_x[2203];
            n_Body_y[2203] = c_Body_y[2203];
            n_Body_x[2204] = c_Body_x[2204];
            n_Body_y[2204] = c_Body_y[2204];
            n_Body_x[2205] = c_Body_x[2205];
            n_Body_y[2205] = c_Body_y[2205];
            n_Body_x[2206] = c_Body_x[2206];
            n_Body_y[2206] = c_Body_y[2206];
            n_Body_x[2207] = c_Body_x[2207];
            n_Body_y[2207] = c_Body_y[2207];
            n_Body_x[2208] = c_Body_x[2208];
            n_Body_y[2208] = c_Body_y[2208];
            n_Body_x[2209] = c_Body_x[2209];
            n_Body_y[2209] = c_Body_y[2209];
            n_Body_x[2210] = c_Body_x[2210];
            n_Body_y[2210] = c_Body_y[2210];
            n_Body_x[2211] = c_Body_x[2211];
            n_Body_y[2211] = c_Body_y[2211];
            n_Body_x[2212] = c_Body_x[2212];
            n_Body_y[2212] = c_Body_y[2212];
            n_Body_x[2213] = c_Body_x[2213];
            n_Body_y[2213] = c_Body_y[2213];
            n_Body_x[2214] = c_Body_x[2214];
            n_Body_y[2214] = c_Body_y[2214];
            n_Body_x[2215] = c_Body_x[2215];
            n_Body_y[2215] = c_Body_y[2215];
            n_Body_x[2216] = c_Body_x[2216];
            n_Body_y[2216] = c_Body_y[2216];
            n_Body_x[2217] = c_Body_x[2217];
            n_Body_y[2217] = c_Body_y[2217];
            n_Body_x[2218] = c_Body_x[2218];
            n_Body_y[2218] = c_Body_y[2218];
            n_Body_x[2219] = c_Body_x[2219];
            n_Body_y[2219] = c_Body_y[2219];
            n_Body_x[2220] = c_Body_x[2220];
            n_Body_y[2220] = c_Body_y[2220];
            n_Body_x[2221] = c_Body_x[2221];
            n_Body_y[2221] = c_Body_y[2221];
            n_Body_x[2222] = c_Body_x[2222];
            n_Body_y[2222] = c_Body_y[2222];
            n_Body_x[2223] = c_Body_x[2223];
            n_Body_y[2223] = c_Body_y[2223];
            n_Body_x[2224] = c_Body_x[2224];
            n_Body_y[2224] = c_Body_y[2224];
            n_Body_x[2225] = c_Body_x[2225];
            n_Body_y[2225] = c_Body_y[2225];
            n_Body_x[2226] = c_Body_x[2226];
            n_Body_y[2226] = c_Body_y[2226];
            n_Body_x[2227] = c_Body_x[2227];
            n_Body_y[2227] = c_Body_y[2227];
            n_Body_x[2228] = c_Body_x[2228];
            n_Body_y[2228] = c_Body_y[2228];
            n_Body_x[2229] = c_Body_x[2229];
            n_Body_y[2229] = c_Body_y[2229];
            n_Body_x[2230] = c_Body_x[2230];
            n_Body_y[2230] = c_Body_y[2230];
            n_Body_x[2231] = c_Body_x[2231];
            n_Body_y[2231] = c_Body_y[2231];
            n_Body_x[2232] = c_Body_x[2232];
            n_Body_y[2232] = c_Body_y[2232];
            n_Body_x[2233] = c_Body_x[2233];
            n_Body_y[2233] = c_Body_y[2233];
            n_Body_x[2234] = c_Body_x[2234];
            n_Body_y[2234] = c_Body_y[2234];
            n_Body_x[2235] = c_Body_x[2235];
            n_Body_y[2235] = c_Body_y[2235];
            n_Body_x[2236] = c_Body_x[2236];
            n_Body_y[2236] = c_Body_y[2236];
            n_Body_x[2237] = c_Body_x[2237];
            n_Body_y[2237] = c_Body_y[2237];
            n_Body_x[2238] = c_Body_x[2238];
            n_Body_y[2238] = c_Body_y[2238];
            n_Body_x[2239] = c_Body_x[2239];
            n_Body_y[2239] = c_Body_y[2239];
            n_Body_x[2240] = c_Body_x[2240];
            n_Body_y[2240] = c_Body_y[2240];
            n_Body_x[2241] = c_Body_x[2241];
            n_Body_y[2241] = c_Body_y[2241];
            n_Body_x[2242] = c_Body_x[2242];
            n_Body_y[2242] = c_Body_y[2242];
            n_Body_x[2243] = c_Body_x[2243];
            n_Body_y[2243] = c_Body_y[2243];
            n_Body_x[2244] = c_Body_x[2244];
            n_Body_y[2244] = c_Body_y[2244];
            n_Body_x[2245] = c_Body_x[2245];
            n_Body_y[2245] = c_Body_y[2245];
            n_Body_x[2246] = c_Body_x[2246];
            n_Body_y[2246] = c_Body_y[2246];
            n_Body_x[2247] = c_Body_x[2247];
            n_Body_y[2247] = c_Body_y[2247];
            n_Body_x[2248] = c_Body_x[2248];
            n_Body_y[2248] = c_Body_y[2248];
            n_Body_x[2249] = c_Body_x[2249];
            n_Body_y[2249] = c_Body_y[2249];
            n_Body_x[2250] = c_Body_x[2250];
            n_Body_y[2250] = c_Body_y[2250];
            n_Body_x[2251] = c_Body_x[2251];
            n_Body_y[2251] = c_Body_y[2251];
            n_Body_x[2252] = c_Body_x[2252];
            n_Body_y[2252] = c_Body_y[2252];
            n_Body_x[2253] = c_Body_x[2253];
            n_Body_y[2253] = c_Body_y[2253];
            n_Body_x[2254] = c_Body_x[2254];
            n_Body_y[2254] = c_Body_y[2254];
            n_Body_x[2255] = c_Body_x[2255];
            n_Body_y[2255] = c_Body_y[2255];
            n_Body_x[2256] = c_Body_x[2256];
            n_Body_y[2256] = c_Body_y[2256];
            n_Body_x[2257] = c_Body_x[2257];
            n_Body_y[2257] = c_Body_y[2257];
            n_Body_x[2258] = c_Body_x[2258];
            n_Body_y[2258] = c_Body_y[2258];
            n_Body_x[2259] = c_Body_x[2259];
            n_Body_y[2259] = c_Body_y[2259];
            n_Body_x[2260] = c_Body_x[2260];
            n_Body_y[2260] = c_Body_y[2260];
            n_Body_x[2261] = c_Body_x[2261];
            n_Body_y[2261] = c_Body_y[2261];
            n_Body_x[2262] = c_Body_x[2262];
            n_Body_y[2262] = c_Body_y[2262];
            n_Body_x[2263] = c_Body_x[2263];
            n_Body_y[2263] = c_Body_y[2263];
            n_Body_x[2264] = c_Body_x[2264];
            n_Body_y[2264] = c_Body_y[2264];
            n_Body_x[2265] = c_Body_x[2265];
            n_Body_y[2265] = c_Body_y[2265];
            n_Body_x[2266] = c_Body_x[2266];
            n_Body_y[2266] = c_Body_y[2266];
            n_Body_x[2267] = c_Body_x[2267];
            n_Body_y[2267] = c_Body_y[2267];
            n_Body_x[2268] = c_Body_x[2268];
            n_Body_y[2268] = c_Body_y[2268];
            n_Body_x[2269] = c_Body_x[2269];
            n_Body_y[2269] = c_Body_y[2269];
            n_Body_x[2270] = c_Body_x[2270];
            n_Body_y[2270] = c_Body_y[2270];
            n_Body_x[2271] = c_Body_x[2271];
            n_Body_y[2271] = c_Body_y[2271];
            n_Body_x[2272] = c_Body_x[2272];
            n_Body_y[2272] = c_Body_y[2272];
            n_Body_x[2273] = c_Body_x[2273];
            n_Body_y[2273] = c_Body_y[2273];
            n_Body_x[2274] = c_Body_x[2274];
            n_Body_y[2274] = c_Body_y[2274];
            n_Body_x[2275] = c_Body_x[2275];
            n_Body_y[2275] = c_Body_y[2275];
            n_Body_x[2276] = c_Body_x[2276];
            n_Body_y[2276] = c_Body_y[2276];
            n_Body_x[2277] = c_Body_x[2277];
            n_Body_y[2277] = c_Body_y[2277];
            n_Body_x[2278] = c_Body_x[2278];
            n_Body_y[2278] = c_Body_y[2278];
            n_Body_x[2279] = c_Body_x[2279];
            n_Body_y[2279] = c_Body_y[2279];
            n_Body_x[2280] = c_Body_x[2280];
            n_Body_y[2280] = c_Body_y[2280];
            n_Body_x[2281] = c_Body_x[2281];
            n_Body_y[2281] = c_Body_y[2281];
            n_Body_x[2282] = c_Body_x[2282];
            n_Body_y[2282] = c_Body_y[2282];
            n_Body_x[2283] = c_Body_x[2283];
            n_Body_y[2283] = c_Body_y[2283];
            n_Body_x[2284] = c_Body_x[2284];
            n_Body_y[2284] = c_Body_y[2284];
            n_Body_x[2285] = c_Body_x[2285];
            n_Body_y[2285] = c_Body_y[2285];
            n_Body_x[2286] = c_Body_x[2286];
            n_Body_y[2286] = c_Body_y[2286];
            n_Body_x[2287] = c_Body_x[2287];
            n_Body_y[2287] = c_Body_y[2287];
            n_Body_x[2288] = c_Body_x[2288];
            n_Body_y[2288] = c_Body_y[2288];
            n_Body_x[2289] = c_Body_x[2289];
            n_Body_y[2289] = c_Body_y[2289];
            n_Body_x[2290] = c_Body_x[2290];
            n_Body_y[2290] = c_Body_y[2290];
            n_Body_x[2291] = c_Body_x[2291];
            n_Body_y[2291] = c_Body_y[2291];
            n_Body_x[2292] = c_Body_x[2292];
            n_Body_y[2292] = c_Body_y[2292];
            n_Body_x[2293] = c_Body_x[2293];
            n_Body_y[2293] = c_Body_y[2293];
            n_Body_x[2294] = c_Body_x[2294];
            n_Body_y[2294] = c_Body_y[2294];
            n_Body_x[2295] = c_Body_x[2295];
            n_Body_y[2295] = c_Body_y[2295];
            n_Body_x[2296] = c_Body_x[2296];
            n_Body_y[2296] = c_Body_y[2296];
            n_Body_x[2297] = c_Body_x[2297];
            n_Body_y[2297] = c_Body_y[2297];
            n_Body_x[2298] = c_Body_x[2298];
            n_Body_y[2298] = c_Body_y[2298];
            n_Body_x[2299] = c_Body_x[2299];
            n_Body_y[2299] = c_Body_y[2299];
            n_Body_x[2300] = c_Body_x[2300];
            n_Body_y[2300] = c_Body_y[2300];
            n_Body_x[2301] = c_Body_x[2301];
            n_Body_y[2301] = c_Body_y[2301];
            n_Body_x[2302] = c_Body_x[2302];
            n_Body_y[2302] = c_Body_y[2302];
            n_Body_x[2303] = c_Body_x[2303];
            n_Body_y[2303] = c_Body_y[2303];
            n_Body_x[2304] = c_Body_x[2304];
            n_Body_y[2304] = c_Body_y[2304];
            n_Body_x[2305] = c_Body_x[2305];
            n_Body_y[2305] = c_Body_y[2305];
            n_Body_x[2306] = c_Body_x[2306];
            n_Body_y[2306] = c_Body_y[2306];
            n_Body_x[2307] = c_Body_x[2307];
            n_Body_y[2307] = c_Body_y[2307];
            n_Body_x[2308] = c_Body_x[2308];
            n_Body_y[2308] = c_Body_y[2308];
            n_Body_x[2309] = c_Body_x[2309];
            n_Body_y[2309] = c_Body_y[2309];
            n_Body_x[2310] = c_Body_x[2310];
            n_Body_y[2310] = c_Body_y[2310];
            n_Body_x[2311] = c_Body_x[2311];
            n_Body_y[2311] = c_Body_y[2311];
            n_Body_x[2312] = c_Body_x[2312];
            n_Body_y[2312] = c_Body_y[2312];
            n_Body_x[2313] = c_Body_x[2313];
            n_Body_y[2313] = c_Body_y[2313];
            n_Body_x[2314] = c_Body_x[2314];
            n_Body_y[2314] = c_Body_y[2314];
            n_Body_x[2315] = c_Body_x[2315];
            n_Body_y[2315] = c_Body_y[2315];
            n_Body_x[2316] = c_Body_x[2316];
            n_Body_y[2316] = c_Body_y[2316];
            n_Body_x[2317] = c_Body_x[2317];
            n_Body_y[2317] = c_Body_y[2317];
            n_Body_x[2318] = c_Body_x[2318];
            n_Body_y[2318] = c_Body_y[2318];
            n_Body_x[2319] = c_Body_x[2319];
            n_Body_y[2319] = c_Body_y[2319];
            n_Body_x[2320] = c_Body_x[2320];
            n_Body_y[2320] = c_Body_y[2320];
            n_Body_x[2321] = c_Body_x[2321];
            n_Body_y[2321] = c_Body_y[2321];
            n_Body_x[2322] = c_Body_x[2322];
            n_Body_y[2322] = c_Body_y[2322];
            n_Body_x[2323] = c_Body_x[2323];
            n_Body_y[2323] = c_Body_y[2323];
            n_Body_x[2324] = c_Body_x[2324];
            n_Body_y[2324] = c_Body_y[2324];
            n_Body_x[2325] = c_Body_x[2325];
            n_Body_y[2325] = c_Body_y[2325];
            n_Body_x[2326] = c_Body_x[2326];
            n_Body_y[2326] = c_Body_y[2326];
            n_Body_x[2327] = c_Body_x[2327];
            n_Body_y[2327] = c_Body_y[2327];
            n_Body_x[2328] = c_Body_x[2328];
            n_Body_y[2328] = c_Body_y[2328];
            n_Body_x[2329] = c_Body_x[2329];
            n_Body_y[2329] = c_Body_y[2329];
            n_Body_x[2330] = c_Body_x[2330];
            n_Body_y[2330] = c_Body_y[2330];
            n_Body_x[2331] = c_Body_x[2331];
            n_Body_y[2331] = c_Body_y[2331];
            n_Body_x[2332] = c_Body_x[2332];
            n_Body_y[2332] = c_Body_y[2332];
            n_Body_x[2333] = c_Body_x[2333];
            n_Body_y[2333] = c_Body_y[2333];
            n_Body_x[2334] = c_Body_x[2334];
            n_Body_y[2334] = c_Body_y[2334];
            n_Body_x[2335] = c_Body_x[2335];
            n_Body_y[2335] = c_Body_y[2335];
            n_Body_x[2336] = c_Body_x[2336];
            n_Body_y[2336] = c_Body_y[2336];
            n_Body_x[2337] = c_Body_x[2337];
            n_Body_y[2337] = c_Body_y[2337];
            n_Body_x[2338] = c_Body_x[2338];
            n_Body_y[2338] = c_Body_y[2338];
            n_Body_x[2339] = c_Body_x[2339];
            n_Body_y[2339] = c_Body_y[2339];
            n_Body_x[2340] = c_Body_x[2340];
            n_Body_y[2340] = c_Body_y[2340];
            n_Body_x[2341] = c_Body_x[2341];
            n_Body_y[2341] = c_Body_y[2341];
            n_Body_x[2342] = c_Body_x[2342];
            n_Body_y[2342] = c_Body_y[2342];
            n_Body_x[2343] = c_Body_x[2343];
            n_Body_y[2343] = c_Body_y[2343];
            n_Body_x[2344] = c_Body_x[2344];
            n_Body_y[2344] = c_Body_y[2344];
            n_Body_x[2345] = c_Body_x[2345];
            n_Body_y[2345] = c_Body_y[2345];
            n_Body_x[2346] = c_Body_x[2346];
            n_Body_y[2346] = c_Body_y[2346];
            n_Body_x[2347] = c_Body_x[2347];
            n_Body_y[2347] = c_Body_y[2347];
            n_Body_x[2348] = c_Body_x[2348];
            n_Body_y[2348] = c_Body_y[2348];
            n_Body_x[2349] = c_Body_x[2349];
            n_Body_y[2349] = c_Body_y[2349];
            n_Body_x[2350] = c_Body_x[2350];
            n_Body_y[2350] = c_Body_y[2350];
            n_Body_x[2351] = c_Body_x[2351];
            n_Body_y[2351] = c_Body_y[2351];
            n_Body_x[2352] = c_Body_x[2352];
            n_Body_y[2352] = c_Body_y[2352];
            n_Body_x[2353] = c_Body_x[2353];
            n_Body_y[2353] = c_Body_y[2353];
            n_Body_x[2354] = c_Body_x[2354];
            n_Body_y[2354] = c_Body_y[2354];
            n_Body_x[2355] = c_Body_x[2355];
            n_Body_y[2355] = c_Body_y[2355];
            n_Body_x[2356] = c_Body_x[2356];
            n_Body_y[2356] = c_Body_y[2356];
            n_Body_x[2357] = c_Body_x[2357];
            n_Body_y[2357] = c_Body_y[2357];
            n_Body_x[2358] = c_Body_x[2358];
            n_Body_y[2358] = c_Body_y[2358];
            n_Body_x[2359] = c_Body_x[2359];
            n_Body_y[2359] = c_Body_y[2359];
            n_Body_x[2360] = c_Body_x[2360];
            n_Body_y[2360] = c_Body_y[2360];
            n_Body_x[2361] = c_Body_x[2361];
            n_Body_y[2361] = c_Body_y[2361];
            n_Body_x[2362] = c_Body_x[2362];
            n_Body_y[2362] = c_Body_y[2362];
            n_Body_x[2363] = c_Body_x[2363];
            n_Body_y[2363] = c_Body_y[2363];
            n_Body_x[2364] = c_Body_x[2364];
            n_Body_y[2364] = c_Body_y[2364];
            n_Body_x[2365] = c_Body_x[2365];
            n_Body_y[2365] = c_Body_y[2365];
            n_Body_x[2366] = c_Body_x[2366];
            n_Body_y[2366] = c_Body_y[2366];
            n_Body_x[2367] = c_Body_x[2367];
            n_Body_y[2367] = c_Body_y[2367];
            n_Body_x[2368] = c_Body_x[2368];
            n_Body_y[2368] = c_Body_y[2368];
            n_Body_x[2369] = c_Body_x[2369];
            n_Body_y[2369] = c_Body_y[2369];
            n_Body_x[2370] = c_Body_x[2370];
            n_Body_y[2370] = c_Body_y[2370];
            n_Body_x[2371] = c_Body_x[2371];
            n_Body_y[2371] = c_Body_y[2371];
            n_Body_x[2372] = c_Body_x[2372];
            n_Body_y[2372] = c_Body_y[2372];
            n_Body_x[2373] = c_Body_x[2373];
            n_Body_y[2373] = c_Body_y[2373];
            n_Body_x[2374] = c_Body_x[2374];
            n_Body_y[2374] = c_Body_y[2374];
            n_Body_x[2375] = c_Body_x[2375];
            n_Body_y[2375] = c_Body_y[2375];
            n_Body_x[2376] = c_Body_x[2376];
            n_Body_y[2376] = c_Body_y[2376];
            n_Body_x[2377] = c_Body_x[2377];
            n_Body_y[2377] = c_Body_y[2377];
            n_Body_x[2378] = c_Body_x[2378];
            n_Body_y[2378] = c_Body_y[2378];
            n_Body_x[2379] = c_Body_x[2379];
            n_Body_y[2379] = c_Body_y[2379];
            n_Body_x[2380] = c_Body_x[2380];
            n_Body_y[2380] = c_Body_y[2380];
            n_Body_x[2381] = c_Body_x[2381];
            n_Body_y[2381] = c_Body_y[2381];
            n_Body_x[2382] = c_Body_x[2382];
            n_Body_y[2382] = c_Body_y[2382];
            n_Body_x[2383] = c_Body_x[2383];
            n_Body_y[2383] = c_Body_y[2383];
            n_Body_x[2384] = c_Body_x[2384];
            n_Body_y[2384] = c_Body_y[2384];
            n_Body_x[2385] = c_Body_x[2385];
            n_Body_y[2385] = c_Body_y[2385];
            n_Body_x[2386] = c_Body_x[2386];
            n_Body_y[2386] = c_Body_y[2386];
            n_Body_x[2387] = c_Body_x[2387];
            n_Body_y[2387] = c_Body_y[2387];
            n_Body_x[2388] = c_Body_x[2388];
            n_Body_y[2388] = c_Body_y[2388];
            n_Body_x[2389] = c_Body_x[2389];
            n_Body_y[2389] = c_Body_y[2389];
            n_Body_x[2390] = c_Body_x[2390];
            n_Body_y[2390] = c_Body_y[2390];
            n_Body_x[2391] = c_Body_x[2391];
            n_Body_y[2391] = c_Body_y[2391];
            n_Body_x[2392] = c_Body_x[2392];
            n_Body_y[2392] = c_Body_y[2392];
            n_Body_x[2393] = c_Body_x[2393];
            n_Body_y[2393] = c_Body_y[2393];
            n_Body_x[2394] = c_Body_x[2394];
            n_Body_y[2394] = c_Body_y[2394];
            n_Body_x[2395] = c_Body_x[2395];
            n_Body_y[2395] = c_Body_y[2395];
            n_Body_x[2396] = c_Body_x[2396];
            n_Body_y[2396] = c_Body_y[2396];
            n_Body_x[2397] = c_Body_x[2397];
            n_Body_y[2397] = c_Body_y[2397];
            n_Body_x[2398] = c_Body_x[2398];
            n_Body_y[2398] = c_Body_y[2398];
            n_Body_x[2399] = c_Body_x[2399];
            n_Body_y[2399] = c_Body_y[2399];
            n_Body_x[2400] = c_Body_x[2400];
            n_Body_y[2400] = c_Body_y[2400];
            n_Body_x[2401] = c_Body_x[2401];
            n_Body_y[2401] = c_Body_y[2401];
            n_Body_x[2402] = c_Body_x[2402];
            n_Body_y[2402] = c_Body_y[2402];
            n_Body_x[2403] = c_Body_x[2403];
            n_Body_y[2403] = c_Body_y[2403];
            n_Body_x[2404] = c_Body_x[2404];
            n_Body_y[2404] = c_Body_y[2404];
            n_Body_x[2405] = c_Body_x[2405];
            n_Body_y[2405] = c_Body_y[2405];
            n_Body_x[2406] = c_Body_x[2406];
            n_Body_y[2406] = c_Body_y[2406];
            n_Body_x[2407] = c_Body_x[2407];
            n_Body_y[2407] = c_Body_y[2407];
            n_Body_x[2408] = c_Body_x[2408];
            n_Body_y[2408] = c_Body_y[2408];
            n_Body_x[2409] = c_Body_x[2409];
            n_Body_y[2409] = c_Body_y[2409];
            n_Body_x[2410] = c_Body_x[2410];
            n_Body_y[2410] = c_Body_y[2410];
            n_Body_x[2411] = c_Body_x[2411];
            n_Body_y[2411] = c_Body_y[2411];
            n_Body_x[2412] = c_Body_x[2412];
            n_Body_y[2412] = c_Body_y[2412];
            n_Body_x[2413] = c_Body_x[2413];
            n_Body_y[2413] = c_Body_y[2413];
            n_Body_x[2414] = c_Body_x[2414];
            n_Body_y[2414] = c_Body_y[2414];
            n_Body_x[2415] = c_Body_x[2415];
            n_Body_y[2415] = c_Body_y[2415];
            n_Body_x[2416] = c_Body_x[2416];
            n_Body_y[2416] = c_Body_y[2416];
            n_Body_x[2417] = c_Body_x[2417];
            n_Body_y[2417] = c_Body_y[2417];
            n_Body_x[2418] = c_Body_x[2418];
            n_Body_y[2418] = c_Body_y[2418];
            n_Body_x[2419] = c_Body_x[2419];
            n_Body_y[2419] = c_Body_y[2419];
            n_Body_x[2420] = c_Body_x[2420];
            n_Body_y[2420] = c_Body_y[2420];
            n_Body_x[2421] = c_Body_x[2421];
            n_Body_y[2421] = c_Body_y[2421];
            n_Body_x[2422] = c_Body_x[2422];
            n_Body_y[2422] = c_Body_y[2422];
            n_Body_x[2423] = c_Body_x[2423];
            n_Body_y[2423] = c_Body_y[2423];
            n_Body_x[2424] = c_Body_x[2424];
            n_Body_y[2424] = c_Body_y[2424];
            n_Body_x[2425] = c_Body_x[2425];
            n_Body_y[2425] = c_Body_y[2425];
            n_Body_x[2426] = c_Body_x[2426];
            n_Body_y[2426] = c_Body_y[2426];
            n_Body_x[2427] = c_Body_x[2427];
            n_Body_y[2427] = c_Body_y[2427];
            n_Body_x[2428] = c_Body_x[2428];
            n_Body_y[2428] = c_Body_y[2428];
            n_Body_x[2429] = c_Body_x[2429];
            n_Body_y[2429] = c_Body_y[2429];
            n_Body_x[2430] = c_Body_x[2430];
            n_Body_y[2430] = c_Body_y[2430];
            n_Body_x[2431] = c_Body_x[2431];
            n_Body_y[2431] = c_Body_y[2431];
            n_Body_x[2432] = c_Body_x[2432];
            n_Body_y[2432] = c_Body_y[2432];
            n_Body_x[2433] = c_Body_x[2433];
            n_Body_y[2433] = c_Body_y[2433];
            n_Body_x[2434] = c_Body_x[2434];
            n_Body_y[2434] = c_Body_y[2434];
            n_Body_x[2435] = c_Body_x[2435];
            n_Body_y[2435] = c_Body_y[2435];
            n_Body_x[2436] = c_Body_x[2436];
            n_Body_y[2436] = c_Body_y[2436];
            n_Body_x[2437] = c_Body_x[2437];
            n_Body_y[2437] = c_Body_y[2437];
            n_Body_x[2438] = c_Body_x[2438];
            n_Body_y[2438] = c_Body_y[2438];
            n_Body_x[2439] = c_Body_x[2439];
            n_Body_y[2439] = c_Body_y[2439];
            n_Body_x[2440] = c_Body_x[2440];
            n_Body_y[2440] = c_Body_y[2440];
            n_Body_x[2441] = c_Body_x[2441];
            n_Body_y[2441] = c_Body_y[2441];
            n_Body_x[2442] = c_Body_x[2442];
            n_Body_y[2442] = c_Body_y[2442];
            n_Body_x[2443] = c_Body_x[2443];
            n_Body_y[2443] = c_Body_y[2443];
            n_Body_x[2444] = c_Body_x[2444];
            n_Body_y[2444] = c_Body_y[2444];
            n_Body_x[2445] = c_Body_x[2445];
            n_Body_y[2445] = c_Body_y[2445];
            n_Body_x[2446] = c_Body_x[2446];
            n_Body_y[2446] = c_Body_y[2446];
            n_Body_x[2447] = c_Body_x[2447];
            n_Body_y[2447] = c_Body_y[2447];
            n_Body_x[2448] = c_Body_x[2448];
            n_Body_y[2448] = c_Body_y[2448];
            n_Body_x[2449] = c_Body_x[2449];
            n_Body_y[2449] = c_Body_y[2449];
            n_Body_x[2450] = c_Body_x[2450];
            n_Body_y[2450] = c_Body_y[2450];
            n_Body_x[2451] = c_Body_x[2451];
            n_Body_y[2451] = c_Body_y[2451];
            n_Body_x[2452] = c_Body_x[2452];
            n_Body_y[2452] = c_Body_y[2452];
            n_Body_x[2453] = c_Body_x[2453];
            n_Body_y[2453] = c_Body_y[2453];
            n_Body_x[2454] = c_Body_x[2454];
            n_Body_y[2454] = c_Body_y[2454];
            n_Body_x[2455] = c_Body_x[2455];
            n_Body_y[2455] = c_Body_y[2455];
            n_Body_x[2456] = c_Body_x[2456];
            n_Body_y[2456] = c_Body_y[2456];
            n_Body_x[2457] = c_Body_x[2457];
            n_Body_y[2457] = c_Body_y[2457];
            n_Body_x[2458] = c_Body_x[2458];
            n_Body_y[2458] = c_Body_y[2458];
            n_Body_x[2459] = c_Body_x[2459];
            n_Body_y[2459] = c_Body_y[2459];
            n_Body_x[2460] = c_Body_x[2460];
            n_Body_y[2460] = c_Body_y[2460];
            n_Body_x[2461] = c_Body_x[2461];
            n_Body_y[2461] = c_Body_y[2461];
            n_Body_x[2462] = c_Body_x[2462];
            n_Body_y[2462] = c_Body_y[2462];
            n_Body_x[2463] = c_Body_x[2463];
            n_Body_y[2463] = c_Body_y[2463];
            n_Body_x[2464] = c_Body_x[2464];
            n_Body_y[2464] = c_Body_y[2464];
            n_Body_x[2465] = c_Body_x[2465];
            n_Body_y[2465] = c_Body_y[2465];
            n_Body_x[2466] = c_Body_x[2466];
            n_Body_y[2466] = c_Body_y[2466];
            n_Body_x[2467] = c_Body_x[2467];
            n_Body_y[2467] = c_Body_y[2467];
            n_Body_x[2468] = c_Body_x[2468];
            n_Body_y[2468] = c_Body_y[2468];
            n_Body_x[2469] = c_Body_x[2469];
            n_Body_y[2469] = c_Body_y[2469];
            n_Body_x[2470] = c_Body_x[2470];
            n_Body_y[2470] = c_Body_y[2470];
            n_Body_x[2471] = c_Body_x[2471];
            n_Body_y[2471] = c_Body_y[2471];
            n_Body_x[2472] = c_Body_x[2472];
            n_Body_y[2472] = c_Body_y[2472];
            n_Body_x[2473] = c_Body_x[2473];
            n_Body_y[2473] = c_Body_y[2473];
            n_Body_x[2474] = c_Body_x[2474];
            n_Body_y[2474] = c_Body_y[2474];
            n_Body_x[2475] = c_Body_x[2475];
            n_Body_y[2475] = c_Body_y[2475];
            n_Body_x[2476] = c_Body_x[2476];
            n_Body_y[2476] = c_Body_y[2476];
            n_Body_x[2477] = c_Body_x[2477];
            n_Body_y[2477] = c_Body_y[2477];
            n_Body_x[2478] = c_Body_x[2478];
            n_Body_y[2478] = c_Body_y[2478];
            n_Body_x[2479] = c_Body_x[2479];
            n_Body_y[2479] = c_Body_y[2479];
            n_Body_x[2480] = c_Body_x[2480];
            n_Body_y[2480] = c_Body_y[2480];
            n_Body_x[2481] = c_Body_x[2481];
            n_Body_y[2481] = c_Body_y[2481];
            n_Body_x[2482] = c_Body_x[2482];
            n_Body_y[2482] = c_Body_y[2482];
            n_Body_x[2483] = c_Body_x[2483];
            n_Body_y[2483] = c_Body_y[2483];
            n_Body_x[2484] = c_Body_x[2484];
            n_Body_y[2484] = c_Body_y[2484];
            n_Body_x[2485] = c_Body_x[2485];
            n_Body_y[2485] = c_Body_y[2485];
            n_Body_x[2486] = c_Body_x[2486];
            n_Body_y[2486] = c_Body_y[2486];
            n_Body_x[2487] = c_Body_x[2487];
            n_Body_y[2487] = c_Body_y[2487];
            n_Body_x[2488] = c_Body_x[2488];
            n_Body_y[2488] = c_Body_y[2488];
            n_Body_x[2489] = c_Body_x[2489];
            n_Body_y[2489] = c_Body_y[2489];
            n_Body_x[2490] = c_Body_x[2490];
            n_Body_y[2490] = c_Body_y[2490];
            n_Body_x[2491] = c_Body_x[2491];
            n_Body_y[2491] = c_Body_y[2491];
            n_Body_x[2492] = c_Body_x[2492];
            n_Body_y[2492] = c_Body_y[2492];
            n_Body_x[2493] = c_Body_x[2493];
            n_Body_y[2493] = c_Body_y[2493];
            n_Body_x[2494] = c_Body_x[2494];
            n_Body_y[2494] = c_Body_y[2494];
            n_Body_x[2495] = c_Body_x[2495];
            n_Body_y[2495] = c_Body_y[2495];
            n_Body_x[2496] = c_Body_x[2496];
            n_Body_y[2496] = c_Body_y[2496];
            n_Body_x[2497] = c_Body_x[2497];
            n_Body_y[2497] = c_Body_y[2497];
            n_Body_x[2498] = c_Body_x[2498];
            n_Body_y[2498] = c_Body_y[2498];
            n_Body_x[2499] = c_Body_x[2499];
            n_Body_y[2499] = c_Body_y[2499];
            n_Body_x[2500] = c_Body_x[2500];
            n_Body_y[2500] = c_Body_y[2500];
            n_Body_x[2501] = c_Body_x[2501];
            n_Body_y[2501] = c_Body_y[2501];
            n_Body_x[2502] = c_Body_x[2502];
            n_Body_y[2502] = c_Body_y[2502];
            n_Body_x[2503] = c_Body_x[2503];
            n_Body_y[2503] = c_Body_y[2503];
            n_Body_x[2504] = c_Body_x[2504];
            n_Body_y[2504] = c_Body_y[2504];
            n_Body_x[2505] = c_Body_x[2505];
            n_Body_y[2505] = c_Body_y[2505];
            n_Body_x[2506] = c_Body_x[2506];
            n_Body_y[2506] = c_Body_y[2506];
            n_Body_x[2507] = c_Body_x[2507];
            n_Body_y[2507] = c_Body_y[2507];
            n_Body_x[2508] = c_Body_x[2508];
            n_Body_y[2508] = c_Body_y[2508];
            n_Body_x[2509] = c_Body_x[2509];
            n_Body_y[2509] = c_Body_y[2509];
            n_Body_x[2510] = c_Body_x[2510];
            n_Body_y[2510] = c_Body_y[2510];
            n_Body_x[2511] = c_Body_x[2511];
            n_Body_y[2511] = c_Body_y[2511];
            n_Body_x[2512] = c_Body_x[2512];
            n_Body_y[2512] = c_Body_y[2512];
            n_Body_x[2513] = c_Body_x[2513];
            n_Body_y[2513] = c_Body_y[2513];
            n_Body_x[2514] = c_Body_x[2514];
            n_Body_y[2514] = c_Body_y[2514];
            n_Body_x[2515] = c_Body_x[2515];
            n_Body_y[2515] = c_Body_y[2515];
            n_Body_x[2516] = c_Body_x[2516];
            n_Body_y[2516] = c_Body_y[2516];
            n_Body_x[2517] = c_Body_x[2517];
            n_Body_y[2517] = c_Body_y[2517];
            n_Body_x[2518] = c_Body_x[2518];
            n_Body_y[2518] = c_Body_y[2518];
            n_Body_x[2519] = c_Body_x[2519];
            n_Body_y[2519] = c_Body_y[2519];
            n_Body_x[2520] = c_Body_x[2520];
            n_Body_y[2520] = c_Body_y[2520];
            n_Body_x[2521] = c_Body_x[2521];
            n_Body_y[2521] = c_Body_y[2521];
            n_Body_x[2522] = c_Body_x[2522];
            n_Body_y[2522] = c_Body_y[2522];
            n_Body_x[2523] = c_Body_x[2523];
            n_Body_y[2523] = c_Body_y[2523];
            n_Body_x[2524] = c_Body_x[2524];
            n_Body_y[2524] = c_Body_y[2524];
            n_Body_x[2525] = c_Body_x[2525];
            n_Body_y[2525] = c_Body_y[2525];
            n_Body_x[2526] = c_Body_x[2526];
            n_Body_y[2526] = c_Body_y[2526];
            n_Body_x[2527] = c_Body_x[2527];
            n_Body_y[2527] = c_Body_y[2527];
            n_Body_x[2528] = c_Body_x[2528];
            n_Body_y[2528] = c_Body_y[2528];
            n_Body_x[2529] = c_Body_x[2529];
            n_Body_y[2529] = c_Body_y[2529];
            n_Body_x[2530] = c_Body_x[2530];
            n_Body_y[2530] = c_Body_y[2530];
            n_Body_x[2531] = c_Body_x[2531];
            n_Body_y[2531] = c_Body_y[2531];
            n_Body_x[2532] = c_Body_x[2532];
            n_Body_y[2532] = c_Body_y[2532];
            n_Body_x[2533] = c_Body_x[2533];
            n_Body_y[2533] = c_Body_y[2533];
            n_Body_x[2534] = c_Body_x[2534];
            n_Body_y[2534] = c_Body_y[2534];
            n_Body_x[2535] = c_Body_x[2535];
            n_Body_y[2535] = c_Body_y[2535];
            n_Body_x[2536] = c_Body_x[2536];
            n_Body_y[2536] = c_Body_y[2536];
            n_Body_x[2537] = c_Body_x[2537];
            n_Body_y[2537] = c_Body_y[2537];
            n_Body_x[2538] = c_Body_x[2538];
            n_Body_y[2538] = c_Body_y[2538];
            n_Body_x[2539] = c_Body_x[2539];
            n_Body_y[2539] = c_Body_y[2539];
            n_Body_x[2540] = c_Body_x[2540];
            n_Body_y[2540] = c_Body_y[2540];
            n_Body_x[2541] = c_Body_x[2541];
            n_Body_y[2541] = c_Body_y[2541];
            n_Body_x[2542] = c_Body_x[2542];
            n_Body_y[2542] = c_Body_y[2542];
            n_Body_x[2543] = c_Body_x[2543];
            n_Body_y[2543] = c_Body_y[2543];
            n_Body_x[2544] = c_Body_x[2544];
            n_Body_y[2544] = c_Body_y[2544];
            n_Body_x[2545] = c_Body_x[2545];
            n_Body_y[2545] = c_Body_y[2545];
            n_Body_x[2546] = c_Body_x[2546];
            n_Body_y[2546] = c_Body_y[2546];
            n_Body_x[2547] = c_Body_x[2547];
            n_Body_y[2547] = c_Body_y[2547];
            n_Body_x[2548] = c_Body_x[2548];
            n_Body_y[2548] = c_Body_y[2548];
            n_Body_x[2549] = c_Body_x[2549];
            n_Body_y[2549] = c_Body_y[2549];
            n_Body_x[2550] = c_Body_x[2550];
            n_Body_y[2550] = c_Body_y[2550];
            n_Body_x[2551] = c_Body_x[2551];
            n_Body_y[2551] = c_Body_y[2551];
            n_Body_x[2552] = c_Body_x[2552];
            n_Body_y[2552] = c_Body_y[2552];
            n_Body_x[2553] = c_Body_x[2553];
            n_Body_y[2553] = c_Body_y[2553];
            n_Body_x[2554] = c_Body_x[2554];
            n_Body_y[2554] = c_Body_y[2554];
            n_Body_x[2555] = c_Body_x[2555];
            n_Body_y[2555] = c_Body_y[2555];
            n_Body_x[2556] = c_Body_x[2556];
            n_Body_y[2556] = c_Body_y[2556];
            n_Body_x[2557] = c_Body_x[2557];
            n_Body_y[2557] = c_Body_y[2557];
            n_Body_x[2558] = c_Body_x[2558];
            n_Body_y[2558] = c_Body_y[2558];
            n_Body_x[2559] = c_Body_x[2559];
            n_Body_y[2559] = c_Body_y[2559];
            n_Body_x[2560] = c_Body_x[2560];
            n_Body_y[2560] = c_Body_y[2560];
            n_Body_x[2561] = c_Body_x[2561];
            n_Body_y[2561] = c_Body_y[2561];
            n_Body_x[2562] = c_Body_x[2562];
            n_Body_y[2562] = c_Body_y[2562];
            n_Body_x[2563] = c_Body_x[2563];
            n_Body_y[2563] = c_Body_y[2563];
            n_Body_x[2564] = c_Body_x[2564];
            n_Body_y[2564] = c_Body_y[2564];
            n_Body_x[2565] = c_Body_x[2565];
            n_Body_y[2565] = c_Body_y[2565];
            n_Body_x[2566] = c_Body_x[2566];
            n_Body_y[2566] = c_Body_y[2566];
            n_Body_x[2567] = c_Body_x[2567];
            n_Body_y[2567] = c_Body_y[2567];
            n_Body_x[2568] = c_Body_x[2568];
            n_Body_y[2568] = c_Body_y[2568];
            n_Body_x[2569] = c_Body_x[2569];
            n_Body_y[2569] = c_Body_y[2569];
            n_Body_x[2570] = c_Body_x[2570];
            n_Body_y[2570] = c_Body_y[2570];
            n_Body_x[2571] = c_Body_x[2571];
            n_Body_y[2571] = c_Body_y[2571];
            n_Body_x[2572] = c_Body_x[2572];
            n_Body_y[2572] = c_Body_y[2572];
            n_Body_x[2573] = c_Body_x[2573];
            n_Body_y[2573] = c_Body_y[2573];
            n_Body_x[2574] = c_Body_x[2574];
            n_Body_y[2574] = c_Body_y[2574];
            n_Body_x[2575] = c_Body_x[2575];
            n_Body_y[2575] = c_Body_y[2575];
            n_Body_x[2576] = c_Body_x[2576];
            n_Body_y[2576] = c_Body_y[2576];
            n_Body_x[2577] = c_Body_x[2577];
            n_Body_y[2577] = c_Body_y[2577];
            n_Body_x[2578] = c_Body_x[2578];
            n_Body_y[2578] = c_Body_y[2578];
            n_Body_x[2579] = c_Body_x[2579];
            n_Body_y[2579] = c_Body_y[2579];
            n_Body_x[2580] = c_Body_x[2580];
            n_Body_y[2580] = c_Body_y[2580];
            n_Body_x[2581] = c_Body_x[2581];
            n_Body_y[2581] = c_Body_y[2581];
            n_Body_x[2582] = c_Body_x[2582];
            n_Body_y[2582] = c_Body_y[2582];
            n_Body_x[2583] = c_Body_x[2583];
            n_Body_y[2583] = c_Body_y[2583];
            n_Body_x[2584] = c_Body_x[2584];
            n_Body_y[2584] = c_Body_y[2584];
            n_Body_x[2585] = c_Body_x[2585];
            n_Body_y[2585] = c_Body_y[2585];
            n_Body_x[2586] = c_Body_x[2586];
            n_Body_y[2586] = c_Body_y[2586];
            n_Body_x[2587] = c_Body_x[2587];
            n_Body_y[2587] = c_Body_y[2587];
            n_Body_x[2588] = c_Body_x[2588];
            n_Body_y[2588] = c_Body_y[2588];
            n_Body_x[2589] = c_Body_x[2589];
            n_Body_y[2589] = c_Body_y[2589];
            n_Body_x[2590] = c_Body_x[2590];
            n_Body_y[2590] = c_Body_y[2590];
            n_Body_x[2591] = c_Body_x[2591];
            n_Body_y[2591] = c_Body_y[2591];
            n_Body_x[2592] = c_Body_x[2592];
            n_Body_y[2592] = c_Body_y[2592];
            n_Body_x[2593] = c_Body_x[2593];
            n_Body_y[2593] = c_Body_y[2593];
            n_Body_x[2594] = c_Body_x[2594];
            n_Body_y[2594] = c_Body_y[2594];
            n_Body_x[2595] = c_Body_x[2595];
            n_Body_y[2595] = c_Body_y[2595];
            n_Body_x[2596] = c_Body_x[2596];
            n_Body_y[2596] = c_Body_y[2596];
            n_Body_x[2597] = c_Body_x[2597];
            n_Body_y[2597] = c_Body_y[2597];
            n_Body_x[2598] = c_Body_x[2598];
            n_Body_y[2598] = c_Body_y[2598];
            n_Body_x[2599] = c_Body_x[2599];
            n_Body_y[2599] = c_Body_y[2599];
            n_Body_x[2600] = c_Body_x[2600];
            n_Body_y[2600] = c_Body_y[2600];
            n_Body_x[2601] = c_Body_x[2601];
            n_Body_y[2601] = c_Body_y[2601];
            n_Body_x[2602] = c_Body_x[2602];
            n_Body_y[2602] = c_Body_y[2602];
            n_Body_x[2603] = c_Body_x[2603];
            n_Body_y[2603] = c_Body_y[2603];
            n_Body_x[2604] = c_Body_x[2604];
            n_Body_y[2604] = c_Body_y[2604];
            n_Body_x[2605] = c_Body_x[2605];
            n_Body_y[2605] = c_Body_y[2605];
            n_Body_x[2606] = c_Body_x[2606];
            n_Body_y[2606] = c_Body_y[2606];
            n_Body_x[2607] = c_Body_x[2607];
            n_Body_y[2607] = c_Body_y[2607];
            n_Body_x[2608] = c_Body_x[2608];
            n_Body_y[2608] = c_Body_y[2608];
            n_Body_x[2609] = c_Body_x[2609];
            n_Body_y[2609] = c_Body_y[2609];
            n_Body_x[2610] = c_Body_x[2610];
            n_Body_y[2610] = c_Body_y[2610];
            n_Body_x[2611] = c_Body_x[2611];
            n_Body_y[2611] = c_Body_y[2611];
            n_Body_x[2612] = c_Body_x[2612];
            n_Body_y[2612] = c_Body_y[2612];
            n_Body_x[2613] = c_Body_x[2613];
            n_Body_y[2613] = c_Body_y[2613];
            n_Body_x[2614] = c_Body_x[2614];
            n_Body_y[2614] = c_Body_y[2614];
            n_Body_x[2615] = c_Body_x[2615];
            n_Body_y[2615] = c_Body_y[2615];
            n_Body_x[2616] = c_Body_x[2616];
            n_Body_y[2616] = c_Body_y[2616];
            n_Body_x[2617] = c_Body_x[2617];
            n_Body_y[2617] = c_Body_y[2617];
            n_Body_x[2618] = c_Body_x[2618];
            n_Body_y[2618] = c_Body_y[2618];
            n_Body_x[2619] = c_Body_x[2619];
            n_Body_y[2619] = c_Body_y[2619];
            n_Body_x[2620] = c_Body_x[2620];
            n_Body_y[2620] = c_Body_y[2620];
            n_Body_x[2621] = c_Body_x[2621];
            n_Body_y[2621] = c_Body_y[2621];
            n_Body_x[2622] = c_Body_x[2622];
            n_Body_y[2622] = c_Body_y[2622];
            n_Body_x[2623] = c_Body_x[2623];
            n_Body_y[2623] = c_Body_y[2623];
            n_Body_x[2624] = c_Body_x[2624];
            n_Body_y[2624] = c_Body_y[2624];
            n_Body_x[2625] = c_Body_x[2625];
            n_Body_y[2625] = c_Body_y[2625];
            n_Body_x[2626] = c_Body_x[2626];
            n_Body_y[2626] = c_Body_y[2626];
            n_Body_x[2627] = c_Body_x[2627];
            n_Body_y[2627] = c_Body_y[2627];
            n_Body_x[2628] = c_Body_x[2628];
            n_Body_y[2628] = c_Body_y[2628];
            n_Body_x[2629] = c_Body_x[2629];
            n_Body_y[2629] = c_Body_y[2629];
            n_Body_x[2630] = c_Body_x[2630];
            n_Body_y[2630] = c_Body_y[2630];
            n_Body_x[2631] = c_Body_x[2631];
            n_Body_y[2631] = c_Body_y[2631];
            n_Body_x[2632] = c_Body_x[2632];
            n_Body_y[2632] = c_Body_y[2632];
            n_Body_x[2633] = c_Body_x[2633];
            n_Body_y[2633] = c_Body_y[2633];
            n_Body_x[2634] = c_Body_x[2634];
            n_Body_y[2634] = c_Body_y[2634];
            n_Body_x[2635] = c_Body_x[2635];
            n_Body_y[2635] = c_Body_y[2635];
            n_Body_x[2636] = c_Body_x[2636];
            n_Body_y[2636] = c_Body_y[2636];
            n_Body_x[2637] = c_Body_x[2637];
            n_Body_y[2637] = c_Body_y[2637];
            n_Body_x[2638] = c_Body_x[2638];
            n_Body_y[2638] = c_Body_y[2638];
            n_Body_x[2639] = c_Body_x[2639];
            n_Body_y[2639] = c_Body_y[2639];
            n_Body_x[2640] = c_Body_x[2640];
            n_Body_y[2640] = c_Body_y[2640];
            n_Body_x[2641] = c_Body_x[2641];
            n_Body_y[2641] = c_Body_y[2641];
            n_Body_x[2642] = c_Body_x[2642];
            n_Body_y[2642] = c_Body_y[2642];
            n_Body_x[2643] = c_Body_x[2643];
            n_Body_y[2643] = c_Body_y[2643];
            n_Body_x[2644] = c_Body_x[2644];
            n_Body_y[2644] = c_Body_y[2644];
            n_Body_x[2645] = c_Body_x[2645];
            n_Body_y[2645] = c_Body_y[2645];
            n_Body_x[2646] = c_Body_x[2646];
            n_Body_y[2646] = c_Body_y[2646];
            n_Body_x[2647] = c_Body_x[2647];
            n_Body_y[2647] = c_Body_y[2647];
            n_Body_x[2648] = c_Body_x[2648];
            n_Body_y[2648] = c_Body_y[2648];
            n_Body_x[2649] = c_Body_x[2649];
            n_Body_y[2649] = c_Body_y[2649];
            n_Body_x[2650] = c_Body_x[2650];
            n_Body_y[2650] = c_Body_y[2650];
            n_Body_x[2651] = c_Body_x[2651];
            n_Body_y[2651] = c_Body_y[2651];
            n_Body_x[2652] = c_Body_x[2652];
            n_Body_y[2652] = c_Body_y[2652];
            n_Body_x[2653] = c_Body_x[2653];
            n_Body_y[2653] = c_Body_y[2653];
            n_Body_x[2654] = c_Body_x[2654];
            n_Body_y[2654] = c_Body_y[2654];
            n_Body_x[2655] = c_Body_x[2655];
            n_Body_y[2655] = c_Body_y[2655];
            n_Body_x[2656] = c_Body_x[2656];
            n_Body_y[2656] = c_Body_y[2656];
            n_Body_x[2657] = c_Body_x[2657];
            n_Body_y[2657] = c_Body_y[2657];
            n_Body_x[2658] = c_Body_x[2658];
            n_Body_y[2658] = c_Body_y[2658];
            n_Body_x[2659] = c_Body_x[2659];
            n_Body_y[2659] = c_Body_y[2659];
            n_Body_x[2660] = c_Body_x[2660];
            n_Body_y[2660] = c_Body_y[2660];
            n_Body_x[2661] = c_Body_x[2661];
            n_Body_y[2661] = c_Body_y[2661];
            n_Body_x[2662] = c_Body_x[2662];
            n_Body_y[2662] = c_Body_y[2662];
            n_Body_x[2663] = c_Body_x[2663];
            n_Body_y[2663] = c_Body_y[2663];
            n_Body_x[2664] = c_Body_x[2664];
            n_Body_y[2664] = c_Body_y[2664];
            n_Body_x[2665] = c_Body_x[2665];
            n_Body_y[2665] = c_Body_y[2665];
            n_Body_x[2666] = c_Body_x[2666];
            n_Body_y[2666] = c_Body_y[2666];
            n_Body_x[2667] = c_Body_x[2667];
            n_Body_y[2667] = c_Body_y[2667];
            n_Body_x[2668] = c_Body_x[2668];
            n_Body_y[2668] = c_Body_y[2668];
            n_Body_x[2669] = c_Body_x[2669];
            n_Body_y[2669] = c_Body_y[2669];
            n_Body_x[2670] = c_Body_x[2670];
            n_Body_y[2670] = c_Body_y[2670];
            n_Body_x[2671] = c_Body_x[2671];
            n_Body_y[2671] = c_Body_y[2671];
            n_Body_x[2672] = c_Body_x[2672];
            n_Body_y[2672] = c_Body_y[2672];
            n_Body_x[2673] = c_Body_x[2673];
            n_Body_y[2673] = c_Body_y[2673];
            n_Body_x[2674] = c_Body_x[2674];
            n_Body_y[2674] = c_Body_y[2674];
            n_Body_x[2675] = c_Body_x[2675];
            n_Body_y[2675] = c_Body_y[2675];
            n_Body_x[2676] = c_Body_x[2676];
            n_Body_y[2676] = c_Body_y[2676];
            n_Body_x[2677] = c_Body_x[2677];
            n_Body_y[2677] = c_Body_y[2677];
            n_Body_x[2678] = c_Body_x[2678];
            n_Body_y[2678] = c_Body_y[2678];
            n_Body_x[2679] = c_Body_x[2679];
            n_Body_y[2679] = c_Body_y[2679];
            n_Body_x[2680] = c_Body_x[2680];
            n_Body_y[2680] = c_Body_y[2680];
            n_Body_x[2681] = c_Body_x[2681];
            n_Body_y[2681] = c_Body_y[2681];
            n_Body_x[2682] = c_Body_x[2682];
            n_Body_y[2682] = c_Body_y[2682];
            n_Body_x[2683] = c_Body_x[2683];
            n_Body_y[2683] = c_Body_y[2683];
            n_Body_x[2684] = c_Body_x[2684];
            n_Body_y[2684] = c_Body_y[2684];
            n_Body_x[2685] = c_Body_x[2685];
            n_Body_y[2685] = c_Body_y[2685];
            n_Body_x[2686] = c_Body_x[2686];
            n_Body_y[2686] = c_Body_y[2686];
            n_Body_x[2687] = c_Body_x[2687];
            n_Body_y[2687] = c_Body_y[2687];
            n_Body_x[2688] = c_Body_x[2688];
            n_Body_y[2688] = c_Body_y[2688];
            n_Body_x[2689] = c_Body_x[2689];
            n_Body_y[2689] = c_Body_y[2689];
            n_Body_x[2690] = c_Body_x[2690];
            n_Body_y[2690] = c_Body_y[2690];
            n_Body_x[2691] = c_Body_x[2691];
            n_Body_y[2691] = c_Body_y[2691];
            n_Body_x[2692] = c_Body_x[2692];
            n_Body_y[2692] = c_Body_y[2692];
            n_Body_x[2693] = c_Body_x[2693];
            n_Body_y[2693] = c_Body_y[2693];
            n_Body_x[2694] = c_Body_x[2694];
            n_Body_y[2694] = c_Body_y[2694];
            n_Body_x[2695] = c_Body_x[2695];
            n_Body_y[2695] = c_Body_y[2695];
            n_Body_x[2696] = c_Body_x[2696];
            n_Body_y[2696] = c_Body_y[2696];
            n_Body_x[2697] = c_Body_x[2697];
            n_Body_y[2697] = c_Body_y[2697];
            n_Body_x[2698] = c_Body_x[2698];
            n_Body_y[2698] = c_Body_y[2698];
            n_Body_x[2699] = c_Body_x[2699];
            n_Body_y[2699] = c_Body_y[2699];
            n_Body_x[2700] = c_Body_x[2700];
            n_Body_y[2700] = c_Body_y[2700];
            n_Body_x[2701] = c_Body_x[2701];
            n_Body_y[2701] = c_Body_y[2701];
            n_Body_x[2702] = c_Body_x[2702];
            n_Body_y[2702] = c_Body_y[2702];
            n_Body_x[2703] = c_Body_x[2703];
            n_Body_y[2703] = c_Body_y[2703];
            n_Body_x[2704] = c_Body_x[2704];
            n_Body_y[2704] = c_Body_y[2704];
            n_Body_x[2705] = c_Body_x[2705];
            n_Body_y[2705] = c_Body_y[2705];
            n_Body_x[2706] = c_Body_x[2706];
            n_Body_y[2706] = c_Body_y[2706];
            n_Body_x[2707] = c_Body_x[2707];
            n_Body_y[2707] = c_Body_y[2707];
            n_Body_x[2708] = c_Body_x[2708];
            n_Body_y[2708] = c_Body_y[2708];
            n_Body_x[2709] = c_Body_x[2709];
            n_Body_y[2709] = c_Body_y[2709];
            n_Body_x[2710] = c_Body_x[2710];
            n_Body_y[2710] = c_Body_y[2710];
            n_Body_x[2711] = c_Body_x[2711];
            n_Body_y[2711] = c_Body_y[2711];
            n_Body_x[2712] = c_Body_x[2712];
            n_Body_y[2712] = c_Body_y[2712];
            n_Body_x[2713] = c_Body_x[2713];
            n_Body_y[2713] = c_Body_y[2713];
            n_Body_x[2714] = c_Body_x[2714];
            n_Body_y[2714] = c_Body_y[2714];
            n_Body_x[2715] = c_Body_x[2715];
            n_Body_y[2715] = c_Body_y[2715];
            n_Body_x[2716] = c_Body_x[2716];
            n_Body_y[2716] = c_Body_y[2716];
            n_Body_x[2717] = c_Body_x[2717];
            n_Body_y[2717] = c_Body_y[2717];
            n_Body_x[2718] = c_Body_x[2718];
            n_Body_y[2718] = c_Body_y[2718];
            n_Body_x[2719] = c_Body_x[2719];
            n_Body_y[2719] = c_Body_y[2719];
            n_Body_x[2720] = c_Body_x[2720];
            n_Body_y[2720] = c_Body_y[2720];
            n_Body_x[2721] = c_Body_x[2721];
            n_Body_y[2721] = c_Body_y[2721];
            n_Body_x[2722] = c_Body_x[2722];
            n_Body_y[2722] = c_Body_y[2722];
            n_Body_x[2723] = c_Body_x[2723];
            n_Body_y[2723] = c_Body_y[2723];
            n_Body_x[2724] = c_Body_x[2724];
            n_Body_y[2724] = c_Body_y[2724];
            n_Body_x[2725] = c_Body_x[2725];
            n_Body_y[2725] = c_Body_y[2725];
            n_Body_x[2726] = c_Body_x[2726];
            n_Body_y[2726] = c_Body_y[2726];
            n_Body_x[2727] = c_Body_x[2727];
            n_Body_y[2727] = c_Body_y[2727];
            n_Body_x[2728] = c_Body_x[2728];
            n_Body_y[2728] = c_Body_y[2728];
            n_Body_x[2729] = c_Body_x[2729];
            n_Body_y[2729] = c_Body_y[2729];
            n_Body_x[2730] = c_Body_x[2730];
            n_Body_y[2730] = c_Body_y[2730];
            n_Body_x[2731] = c_Body_x[2731];
            n_Body_y[2731] = c_Body_y[2731];
            n_Body_x[2732] = c_Body_x[2732];
            n_Body_y[2732] = c_Body_y[2732];
            n_Body_x[2733] = c_Body_x[2733];
            n_Body_y[2733] = c_Body_y[2733];
            n_Body_x[2734] = c_Body_x[2734];
            n_Body_y[2734] = c_Body_y[2734];
            n_Body_x[2735] = c_Body_x[2735];
            n_Body_y[2735] = c_Body_y[2735];
            n_Body_x[2736] = c_Body_x[2736];
            n_Body_y[2736] = c_Body_y[2736];
            n_Body_x[2737] = c_Body_x[2737];
            n_Body_y[2737] = c_Body_y[2737];
            n_Body_x[2738] = c_Body_x[2738];
            n_Body_y[2738] = c_Body_y[2738];
            n_Body_x[2739] = c_Body_x[2739];
            n_Body_y[2739] = c_Body_y[2739];
            n_Body_x[2740] = c_Body_x[2740];
            n_Body_y[2740] = c_Body_y[2740];
            n_Body_x[2741] = c_Body_x[2741];
            n_Body_y[2741] = c_Body_y[2741];
            n_Body_x[2742] = c_Body_x[2742];
            n_Body_y[2742] = c_Body_y[2742];
            n_Body_x[2743] = c_Body_x[2743];
            n_Body_y[2743] = c_Body_y[2743];
            n_Body_x[2744] = c_Body_x[2744];
            n_Body_y[2744] = c_Body_y[2744];
            n_Body_x[2745] = c_Body_x[2745];
            n_Body_y[2745] = c_Body_y[2745];
            n_Body_x[2746] = c_Body_x[2746];
            n_Body_y[2746] = c_Body_y[2746];
            n_Body_x[2747] = c_Body_x[2747];
            n_Body_y[2747] = c_Body_y[2747];
            n_Body_x[2748] = c_Body_x[2748];
            n_Body_y[2748] = c_Body_y[2748];
            n_Body_x[2749] = c_Body_x[2749];
            n_Body_y[2749] = c_Body_y[2749];
            n_Body_x[2750] = c_Body_x[2750];
            n_Body_y[2750] = c_Body_y[2750];
            n_Body_x[2751] = c_Body_x[2751];
            n_Body_y[2751] = c_Body_y[2751];
            n_Body_x[2752] = c_Body_x[2752];
            n_Body_y[2752] = c_Body_y[2752];
            n_Body_x[2753] = c_Body_x[2753];
            n_Body_y[2753] = c_Body_y[2753];
            n_Body_x[2754] = c_Body_x[2754];
            n_Body_y[2754] = c_Body_y[2754];
            n_Body_x[2755] = c_Body_x[2755];
            n_Body_y[2755] = c_Body_y[2755];
            n_Body_x[2756] = c_Body_x[2756];
            n_Body_y[2756] = c_Body_y[2756];
            n_Body_x[2757] = c_Body_x[2757];
            n_Body_y[2757] = c_Body_y[2757];
            n_Body_x[2758] = c_Body_x[2758];
            n_Body_y[2758] = c_Body_y[2758];
            n_Body_x[2759] = c_Body_x[2759];
            n_Body_y[2759] = c_Body_y[2759];
            n_Body_x[2760] = c_Body_x[2760];
            n_Body_y[2760] = c_Body_y[2760];
            n_Body_x[2761] = c_Body_x[2761];
            n_Body_y[2761] = c_Body_y[2761];
            n_Body_x[2762] = c_Body_x[2762];
            n_Body_y[2762] = c_Body_y[2762];
            n_Body_x[2763] = c_Body_x[2763];
            n_Body_y[2763] = c_Body_y[2763];
            n_Body_x[2764] = c_Body_x[2764];
            n_Body_y[2764] = c_Body_y[2764];
            n_Body_x[2765] = c_Body_x[2765];
            n_Body_y[2765] = c_Body_y[2765];
            n_Body_x[2766] = c_Body_x[2766];
            n_Body_y[2766] = c_Body_y[2766];
            n_Body_x[2767] = c_Body_x[2767];
            n_Body_y[2767] = c_Body_y[2767];
            n_Body_x[2768] = c_Body_x[2768];
            n_Body_y[2768] = c_Body_y[2768];
            n_Body_x[2769] = c_Body_x[2769];
            n_Body_y[2769] = c_Body_y[2769];
            n_Body_x[2770] = c_Body_x[2770];
            n_Body_y[2770] = c_Body_y[2770];
            n_Body_x[2771] = c_Body_x[2771];
            n_Body_y[2771] = c_Body_y[2771];
            n_Body_x[2772] = c_Body_x[2772];
            n_Body_y[2772] = c_Body_y[2772];
            n_Body_x[2773] = c_Body_x[2773];
            n_Body_y[2773] = c_Body_y[2773];
            n_Body_x[2774] = c_Body_x[2774];
            n_Body_y[2774] = c_Body_y[2774];
            n_Body_x[2775] = c_Body_x[2775];
            n_Body_y[2775] = c_Body_y[2775];
            n_Body_x[2776] = c_Body_x[2776];
            n_Body_y[2776] = c_Body_y[2776];
            n_Body_x[2777] = c_Body_x[2777];
            n_Body_y[2777] = c_Body_y[2777];
            n_Body_x[2778] = c_Body_x[2778];
            n_Body_y[2778] = c_Body_y[2778];
            n_Body_x[2779] = c_Body_x[2779];
            n_Body_y[2779] = c_Body_y[2779];
            n_Body_x[2780] = c_Body_x[2780];
            n_Body_y[2780] = c_Body_y[2780];
            n_Body_x[2781] = c_Body_x[2781];
            n_Body_y[2781] = c_Body_y[2781];
            n_Body_x[2782] = c_Body_x[2782];
            n_Body_y[2782] = c_Body_y[2782];
            n_Body_x[2783] = c_Body_x[2783];
            n_Body_y[2783] = c_Body_y[2783];
            n_Body_x[2784] = c_Body_x[2784];
            n_Body_y[2784] = c_Body_y[2784];
            n_Body_x[2785] = c_Body_x[2785];
            n_Body_y[2785] = c_Body_y[2785];
            n_Body_x[2786] = c_Body_x[2786];
            n_Body_y[2786] = c_Body_y[2786];
            n_Body_x[2787] = c_Body_x[2787];
            n_Body_y[2787] = c_Body_y[2787];
            n_Body_x[2788] = c_Body_x[2788];
            n_Body_y[2788] = c_Body_y[2788];
            n_Body_x[2789] = c_Body_x[2789];
            n_Body_y[2789] = c_Body_y[2789];
            n_Body_x[2790] = c_Body_x[2790];
            n_Body_y[2790] = c_Body_y[2790];
            n_Body_x[2791] = c_Body_x[2791];
            n_Body_y[2791] = c_Body_y[2791];
            n_Body_x[2792] = c_Body_x[2792];
            n_Body_y[2792] = c_Body_y[2792];
            n_Body_x[2793] = c_Body_x[2793];
            n_Body_y[2793] = c_Body_y[2793];
            n_Body_x[2794] = c_Body_x[2794];
            n_Body_y[2794] = c_Body_y[2794];
            n_Body_x[2795] = c_Body_x[2795];
            n_Body_y[2795] = c_Body_y[2795];
            n_Body_x[2796] = c_Body_x[2796];
            n_Body_y[2796] = c_Body_y[2796];
            n_Body_x[2797] = c_Body_x[2797];
            n_Body_y[2797] = c_Body_y[2797];
            n_Body_x[2798] = c_Body_x[2798];
            n_Body_y[2798] = c_Body_y[2798];
            n_Body_x[2799] = c_Body_x[2799];
            n_Body_y[2799] = c_Body_y[2799];
            n_Body_x[2800] = c_Body_x[2800];
            n_Body_y[2800] = c_Body_y[2800];
            n_Body_x[2801] = c_Body_x[2801];
            n_Body_y[2801] = c_Body_y[2801];
            n_Body_x[2802] = c_Body_x[2802];
            n_Body_y[2802] = c_Body_y[2802];
            n_Body_x[2803] = c_Body_x[2803];
            n_Body_y[2803] = c_Body_y[2803];
            n_Body_x[2804] = c_Body_x[2804];
            n_Body_y[2804] = c_Body_y[2804];
            n_Body_x[2805] = c_Body_x[2805];
            n_Body_y[2805] = c_Body_y[2805];
            n_Body_x[2806] = c_Body_x[2806];
            n_Body_y[2806] = c_Body_y[2806];
            n_Body_x[2807] = c_Body_x[2807];
            n_Body_y[2807] = c_Body_y[2807];
            n_Body_x[2808] = c_Body_x[2808];
            n_Body_y[2808] = c_Body_y[2808];
            n_Body_x[2809] = c_Body_x[2809];
            n_Body_y[2809] = c_Body_y[2809];
            n_Body_x[2810] = c_Body_x[2810];
            n_Body_y[2810] = c_Body_y[2810];
            n_Body_x[2811] = c_Body_x[2811];
            n_Body_y[2811] = c_Body_y[2811];
            n_Body_x[2812] = c_Body_x[2812];
            n_Body_y[2812] = c_Body_y[2812];
            n_Body_x[2813] = c_Body_x[2813];
            n_Body_y[2813] = c_Body_y[2813];
            n_Body_x[2814] = c_Body_x[2814];
            n_Body_y[2814] = c_Body_y[2814];
            n_Body_x[2815] = c_Body_x[2815];
            n_Body_y[2815] = c_Body_y[2815];
            n_Body_x[2816] = c_Body_x[2816];
            n_Body_y[2816] = c_Body_y[2816];
            n_Body_x[2817] = c_Body_x[2817];
            n_Body_y[2817] = c_Body_y[2817];
            n_Body_x[2818] = c_Body_x[2818];
            n_Body_y[2818] = c_Body_y[2818];
            n_Body_x[2819] = c_Body_x[2819];
            n_Body_y[2819] = c_Body_y[2819];
            n_Body_x[2820] = c_Body_x[2820];
            n_Body_y[2820] = c_Body_y[2820];
            n_Body_x[2821] = c_Body_x[2821];
            n_Body_y[2821] = c_Body_y[2821];
            n_Body_x[2822] = c_Body_x[2822];
            n_Body_y[2822] = c_Body_y[2822];
            n_Body_x[2823] = c_Body_x[2823];
            n_Body_y[2823] = c_Body_y[2823];
            n_Body_x[2824] = c_Body_x[2824];
            n_Body_y[2824] = c_Body_y[2824];
            n_Body_x[2825] = c_Body_x[2825];
            n_Body_y[2825] = c_Body_y[2825];
            n_Body_x[2826] = c_Body_x[2826];
            n_Body_y[2826] = c_Body_y[2826];
            n_Body_x[2827] = c_Body_x[2827];
            n_Body_y[2827] = c_Body_y[2827];
            n_Body_x[2828] = c_Body_x[2828];
            n_Body_y[2828] = c_Body_y[2828];
            n_Body_x[2829] = c_Body_x[2829];
            n_Body_y[2829] = c_Body_y[2829];
            n_Body_x[2830] = c_Body_x[2830];
            n_Body_y[2830] = c_Body_y[2830];
            n_Body_x[2831] = c_Body_x[2831];
            n_Body_y[2831] = c_Body_y[2831];
            n_Body_x[2832] = c_Body_x[2832];
            n_Body_y[2832] = c_Body_y[2832];
            n_Body_x[2833] = c_Body_x[2833];
            n_Body_y[2833] = c_Body_y[2833];
            n_Body_x[2834] = c_Body_x[2834];
            n_Body_y[2834] = c_Body_y[2834];
            n_Body_x[2835] = c_Body_x[2835];
            n_Body_y[2835] = c_Body_y[2835];
            n_Body_x[2836] = c_Body_x[2836];
            n_Body_y[2836] = c_Body_y[2836];
            n_Body_x[2837] = c_Body_x[2837];
            n_Body_y[2837] = c_Body_y[2837];
            n_Body_x[2838] = c_Body_x[2838];
            n_Body_y[2838] = c_Body_y[2838];
            n_Body_x[2839] = c_Body_x[2839];
            n_Body_y[2839] = c_Body_y[2839];
            n_Body_x[2840] = c_Body_x[2840];
            n_Body_y[2840] = c_Body_y[2840];
            n_Body_x[2841] = c_Body_x[2841];
            n_Body_y[2841] = c_Body_y[2841];
            n_Body_x[2842] = c_Body_x[2842];
            n_Body_y[2842] = c_Body_y[2842];
            n_Body_x[2843] = c_Body_x[2843];
            n_Body_y[2843] = c_Body_y[2843];
            n_Body_x[2844] = c_Body_x[2844];
            n_Body_y[2844] = c_Body_y[2844];
            n_Body_x[2845] = c_Body_x[2845];
            n_Body_y[2845] = c_Body_y[2845];
            n_Body_x[2846] = c_Body_x[2846];
            n_Body_y[2846] = c_Body_y[2846];
            n_Body_x[2847] = c_Body_x[2847];
            n_Body_y[2847] = c_Body_y[2847];
            n_Body_x[2848] = c_Body_x[2848];
            n_Body_y[2848] = c_Body_y[2848];
            n_Body_x[2849] = c_Body_x[2849];
            n_Body_y[2849] = c_Body_y[2849];
            n_Body_x[2850] = c_Body_x[2850];
            n_Body_y[2850] = c_Body_y[2850];
            n_Body_x[2851] = c_Body_x[2851];
            n_Body_y[2851] = c_Body_y[2851];
            n_Body_x[2852] = c_Body_x[2852];
            n_Body_y[2852] = c_Body_y[2852];
            n_Body_x[2853] = c_Body_x[2853];
            n_Body_y[2853] = c_Body_y[2853];
            n_Body_x[2854] = c_Body_x[2854];
            n_Body_y[2854] = c_Body_y[2854];
            n_Body_x[2855] = c_Body_x[2855];
            n_Body_y[2855] = c_Body_y[2855];
            n_Body_x[2856] = c_Body_x[2856];
            n_Body_y[2856] = c_Body_y[2856];
            n_Body_x[2857] = c_Body_x[2857];
            n_Body_y[2857] = c_Body_y[2857];
            n_Body_x[2858] = c_Body_x[2858];
            n_Body_y[2858] = c_Body_y[2858];
            n_Body_x[2859] = c_Body_x[2859];
            n_Body_y[2859] = c_Body_y[2859];
            n_Body_x[2860] = c_Body_x[2860];
            n_Body_y[2860] = c_Body_y[2860];
            n_Body_x[2861] = c_Body_x[2861];
            n_Body_y[2861] = c_Body_y[2861];
            n_Body_x[2862] = c_Body_x[2862];
            n_Body_y[2862] = c_Body_y[2862];
            n_Body_x[2863] = c_Body_x[2863];
            n_Body_y[2863] = c_Body_y[2863];
            n_Body_x[2864] = c_Body_x[2864];
            n_Body_y[2864] = c_Body_y[2864];
            n_Body_x[2865] = c_Body_x[2865];
            n_Body_y[2865] = c_Body_y[2865];
            n_Body_x[2866] = c_Body_x[2866];
            n_Body_y[2866] = c_Body_y[2866];
            n_Body_x[2867] = c_Body_x[2867];
            n_Body_y[2867] = c_Body_y[2867];
            n_Body_x[2868] = c_Body_x[2868];
            n_Body_y[2868] = c_Body_y[2868];
            n_Body_x[2869] = c_Body_x[2869];
            n_Body_y[2869] = c_Body_y[2869];
            n_Body_x[2870] = c_Body_x[2870];
            n_Body_y[2870] = c_Body_y[2870];
            n_Body_x[2871] = c_Body_x[2871];
            n_Body_y[2871] = c_Body_y[2871];
            n_Body_x[2872] = c_Body_x[2872];
            n_Body_y[2872] = c_Body_y[2872];
            n_Body_x[2873] = c_Body_x[2873];
            n_Body_y[2873] = c_Body_y[2873];
            n_Body_x[2874] = c_Body_x[2874];
            n_Body_y[2874] = c_Body_y[2874];
            n_Body_x[2875] = c_Body_x[2875];
            n_Body_y[2875] = c_Body_y[2875];
            n_Body_x[2876] = c_Body_x[2876];
            n_Body_y[2876] = c_Body_y[2876];
            n_Body_x[2877] = c_Body_x[2877];
            n_Body_y[2877] = c_Body_y[2877];
            n_Body_x[2878] = c_Body_x[2878];
            n_Body_y[2878] = c_Body_y[2878];
            n_Body_x[2879] = c_Body_x[2879];
            n_Body_y[2879] = c_Body_y[2879];
            n_Body_x[2880] = c_Body_x[2880];
            n_Body_y[2880] = c_Body_y[2880];
            n_Body_x[2881] = c_Body_x[2881];
            n_Body_y[2881] = c_Body_y[2881];
            n_Body_x[2882] = c_Body_x[2882];
            n_Body_y[2882] = c_Body_y[2882];
            n_Body_x[2883] = c_Body_x[2883];
            n_Body_y[2883] = c_Body_y[2883];
            n_Body_x[2884] = c_Body_x[2884];
            n_Body_y[2884] = c_Body_y[2884];
            n_Body_x[2885] = c_Body_x[2885];
            n_Body_y[2885] = c_Body_y[2885];
            n_Body_x[2886] = c_Body_x[2886];
            n_Body_y[2886] = c_Body_y[2886];
            n_Body_x[2887] = c_Body_x[2887];
            n_Body_y[2887] = c_Body_y[2887];
            n_Body_x[2888] = c_Body_x[2888];
            n_Body_y[2888] = c_Body_y[2888];
            n_Body_x[2889] = c_Body_x[2889];
            n_Body_y[2889] = c_Body_y[2889];
            n_Body_x[2890] = c_Body_x[2890];
            n_Body_y[2890] = c_Body_y[2890];
            n_Body_x[2891] = c_Body_x[2891];
            n_Body_y[2891] = c_Body_y[2891];
            n_Body_x[2892] = c_Body_x[2892];
            n_Body_y[2892] = c_Body_y[2892];
            n_Body_x[2893] = c_Body_x[2893];
            n_Body_y[2893] = c_Body_y[2893];
            n_Body_x[2894] = c_Body_x[2894];
            n_Body_y[2894] = c_Body_y[2894];
            n_Body_x[2895] = c_Body_x[2895];
            n_Body_y[2895] = c_Body_y[2895];
            n_Body_x[2896] = c_Body_x[2896];
            n_Body_y[2896] = c_Body_y[2896];
            n_Body_x[2897] = c_Body_x[2897];
            n_Body_y[2897] = c_Body_y[2897];
            n_Body_x[2898] = c_Body_x[2898];
            n_Body_y[2898] = c_Body_y[2898];
            n_Body_x[2899] = c_Body_x[2899];
            n_Body_y[2899] = c_Body_y[2899];
            n_Body_x[2900] = c_Body_x[2900];
            n_Body_y[2900] = c_Body_y[2900];
            n_Body_x[2901] = c_Body_x[2901];
            n_Body_y[2901] = c_Body_y[2901];
            n_Body_x[2902] = c_Body_x[2902];
            n_Body_y[2902] = c_Body_y[2902];
            n_Body_x[2903] = c_Body_x[2903];
            n_Body_y[2903] = c_Body_y[2903];
            n_Body_x[2904] = c_Body_x[2904];
            n_Body_y[2904] = c_Body_y[2904];
            n_Body_x[2905] = c_Body_x[2905];
            n_Body_y[2905] = c_Body_y[2905];
            n_Body_x[2906] = c_Body_x[2906];
            n_Body_y[2906] = c_Body_y[2906];
            n_Body_x[2907] = c_Body_x[2907];
            n_Body_y[2907] = c_Body_y[2907];
            n_Body_x[2908] = c_Body_x[2908];
            n_Body_y[2908] = c_Body_y[2908];
            n_Body_x[2909] = c_Body_x[2909];
            n_Body_y[2909] = c_Body_y[2909];
            n_Body_x[2910] = c_Body_x[2910];
            n_Body_y[2910] = c_Body_y[2910];
            n_Body_x[2911] = c_Body_x[2911];
            n_Body_y[2911] = c_Body_y[2911];
            n_Body_x[2912] = c_Body_x[2912];
            n_Body_y[2912] = c_Body_y[2912];
            n_Body_x[2913] = c_Body_x[2913];
            n_Body_y[2913] = c_Body_y[2913];
            n_Body_x[2914] = c_Body_x[2914];
            n_Body_y[2914] = c_Body_y[2914];
            n_Body_x[2915] = c_Body_x[2915];
            n_Body_y[2915] = c_Body_y[2915];
            n_Body_x[2916] = c_Body_x[2916];
            n_Body_y[2916] = c_Body_y[2916];
            n_Body_x[2917] = c_Body_x[2917];
            n_Body_y[2917] = c_Body_y[2917];
            n_Body_x[2918] = c_Body_x[2918];
            n_Body_y[2918] = c_Body_y[2918];
            n_Body_x[2919] = c_Body_x[2919];
            n_Body_y[2919] = c_Body_y[2919];
            n_Body_x[2920] = c_Body_x[2920];
            n_Body_y[2920] = c_Body_y[2920];
            n_Body_x[2921] = c_Body_x[2921];
            n_Body_y[2921] = c_Body_y[2921];
            n_Body_x[2922] = c_Body_x[2922];
            n_Body_y[2922] = c_Body_y[2922];
            n_Body_x[2923] = c_Body_x[2923];
            n_Body_y[2923] = c_Body_y[2923];
            n_Body_x[2924] = c_Body_x[2924];
            n_Body_y[2924] = c_Body_y[2924];
            n_Body_x[2925] = c_Body_x[2925];
            n_Body_y[2925] = c_Body_y[2925];
            n_Body_x[2926] = c_Body_x[2926];
            n_Body_y[2926] = c_Body_y[2926];
            n_Body_x[2927] = c_Body_x[2927];
            n_Body_y[2927] = c_Body_y[2927];
            n_Body_x[2928] = c_Body_x[2928];
            n_Body_y[2928] = c_Body_y[2928];
            n_Body_x[2929] = c_Body_x[2929];
            n_Body_y[2929] = c_Body_y[2929];
            n_Body_x[2930] = c_Body_x[2930];
            n_Body_y[2930] = c_Body_y[2930];
            n_Body_x[2931] = c_Body_x[2931];
            n_Body_y[2931] = c_Body_y[2931];
            n_Body_x[2932] = c_Body_x[2932];
            n_Body_y[2932] = c_Body_y[2932];
            n_Body_x[2933] = c_Body_x[2933];
            n_Body_y[2933] = c_Body_y[2933];
            n_Body_x[2934] = c_Body_x[2934];
            n_Body_y[2934] = c_Body_y[2934];
            n_Body_x[2935] = c_Body_x[2935];
            n_Body_y[2935] = c_Body_y[2935];
            n_Body_x[2936] = c_Body_x[2936];
            n_Body_y[2936] = c_Body_y[2936];
            n_Body_x[2937] = c_Body_x[2937];
            n_Body_y[2937] = c_Body_y[2937];
            n_Body_x[2938] = c_Body_x[2938];
            n_Body_y[2938] = c_Body_y[2938];
            n_Body_x[2939] = c_Body_x[2939];
            n_Body_y[2939] = c_Body_y[2939];
            n_Body_x[2940] = c_Body_x[2940];
            n_Body_y[2940] = c_Body_y[2940];
            n_Body_x[2941] = c_Body_x[2941];
            n_Body_y[2941] = c_Body_y[2941];
            n_Body_x[2942] = c_Body_x[2942];
            n_Body_y[2942] = c_Body_y[2942];
            n_Body_x[2943] = c_Body_x[2943];
            n_Body_y[2943] = c_Body_y[2943];
            n_Body_x[2944] = c_Body_x[2944];
            n_Body_y[2944] = c_Body_y[2944];
            n_Body_x[2945] = c_Body_x[2945];
            n_Body_y[2945] = c_Body_y[2945];
            n_Body_x[2946] = c_Body_x[2946];
            n_Body_y[2946] = c_Body_y[2946];
            n_Body_x[2947] = c_Body_x[2947];
            n_Body_y[2947] = c_Body_y[2947];
            n_Body_x[2948] = c_Body_x[2948];
            n_Body_y[2948] = c_Body_y[2948];
            n_Body_x[2949] = c_Body_x[2949];
            n_Body_y[2949] = c_Body_y[2949];
            n_Body_x[2950] = c_Body_x[2950];
            n_Body_y[2950] = c_Body_y[2950];
            n_Body_x[2951] = c_Body_x[2951];
            n_Body_y[2951] = c_Body_y[2951];
            n_Body_x[2952] = c_Body_x[2952];
            n_Body_y[2952] = c_Body_y[2952];
            n_Body_x[2953] = c_Body_x[2953];
            n_Body_y[2953] = c_Body_y[2953];
            n_Body_x[2954] = c_Body_x[2954];
            n_Body_y[2954] = c_Body_y[2954];
            n_Body_x[2955] = c_Body_x[2955];
            n_Body_y[2955] = c_Body_y[2955];
            n_Body_x[2956] = c_Body_x[2956];
            n_Body_y[2956] = c_Body_y[2956];
            n_Body_x[2957] = c_Body_x[2957];
            n_Body_y[2957] = c_Body_y[2957];
            n_Body_x[2958] = c_Body_x[2958];
            n_Body_y[2958] = c_Body_y[2958];
            n_Body_x[2959] = c_Body_x[2959];
            n_Body_y[2959] = c_Body_y[2959];
            n_Body_x[2960] = c_Body_x[2960];
            n_Body_y[2960] = c_Body_y[2960];
            n_Body_x[2961] = c_Body_x[2961];
            n_Body_y[2961] = c_Body_y[2961];
            n_Body_x[2962] = c_Body_x[2962];
            n_Body_y[2962] = c_Body_y[2962];
            n_Body_x[2963] = c_Body_x[2963];
            n_Body_y[2963] = c_Body_y[2963];
            n_Body_x[2964] = c_Body_x[2964];
            n_Body_y[2964] = c_Body_y[2964];
            n_Body_x[2965] = c_Body_x[2965];
            n_Body_y[2965] = c_Body_y[2965];
            n_Body_x[2966] = c_Body_x[2966];
            n_Body_y[2966] = c_Body_y[2966];
            n_Body_x[2967] = c_Body_x[2967];
            n_Body_y[2967] = c_Body_y[2967];
            n_Body_x[2968] = c_Body_x[2968];
            n_Body_y[2968] = c_Body_y[2968];
            n_Body_x[2969] = c_Body_x[2969];
            n_Body_y[2969] = c_Body_y[2969];
            n_Body_x[2970] = c_Body_x[2970];
            n_Body_y[2970] = c_Body_y[2970];
            n_Body_x[2971] = c_Body_x[2971];
            n_Body_y[2971] = c_Body_y[2971];
            n_Body_x[2972] = c_Body_x[2972];
            n_Body_y[2972] = c_Body_y[2972];
            n_Body_x[2973] = c_Body_x[2973];
            n_Body_y[2973] = c_Body_y[2973];
            n_Body_x[2974] = c_Body_x[2974];
            n_Body_y[2974] = c_Body_y[2974];
            n_Body_x[2975] = c_Body_x[2975];
            n_Body_y[2975] = c_Body_y[2975];
            n_Body_x[2976] = c_Body_x[2976];
            n_Body_y[2976] = c_Body_y[2976];
            n_Body_x[2977] = c_Body_x[2977];
            n_Body_y[2977] = c_Body_y[2977];
            n_Body_x[2978] = c_Body_x[2978];
            n_Body_y[2978] = c_Body_y[2978];
            n_Body_x[2979] = c_Body_x[2979];
            n_Body_y[2979] = c_Body_y[2979];
            n_Body_x[2980] = c_Body_x[2980];
            n_Body_y[2980] = c_Body_y[2980];
            n_Body_x[2981] = c_Body_x[2981];
            n_Body_y[2981] = c_Body_y[2981];
            n_Body_x[2982] = c_Body_x[2982];
            n_Body_y[2982] = c_Body_y[2982];
            n_Body_x[2983] = c_Body_x[2983];
            n_Body_y[2983] = c_Body_y[2983];
            n_Body_x[2984] = c_Body_x[2984];
            n_Body_y[2984] = c_Body_y[2984];
            n_Body_x[2985] = c_Body_x[2985];
            n_Body_y[2985] = c_Body_y[2985];
            n_Body_x[2986] = c_Body_x[2986];
            n_Body_y[2986] = c_Body_y[2986];
            n_Body_x[2987] = c_Body_x[2987];
            n_Body_y[2987] = c_Body_y[2987];
            n_Body_x[2988] = c_Body_x[2988];
            n_Body_y[2988] = c_Body_y[2988];
            n_Body_x[2989] = c_Body_x[2989];
            n_Body_y[2989] = c_Body_y[2989];
            n_Body_x[2990] = c_Body_x[2990];
            n_Body_y[2990] = c_Body_y[2990];
            n_Body_x[2991] = c_Body_x[2991];
            n_Body_y[2991] = c_Body_y[2991];
            n_Body_x[2992] = c_Body_x[2992];
            n_Body_y[2992] = c_Body_y[2992];
            n_Body_x[2993] = c_Body_x[2993];
            n_Body_y[2993] = c_Body_y[2993];
            n_Body_x[2994] = c_Body_x[2994];
            n_Body_y[2994] = c_Body_y[2994];
            n_Body_x[2995] = c_Body_x[2995];
            n_Body_y[2995] = c_Body_y[2995];
            n_Body_x[2996] = c_Body_x[2996];
            n_Body_y[2996] = c_Body_y[2996];
            n_Body_x[2997] = c_Body_x[2997];
            n_Body_y[2997] = c_Body_y[2997];
            n_Body_x[2998] = c_Body_x[2998];
            n_Body_y[2998] = c_Body_y[2998];
            n_Body_x[2999] = c_Body_x[2999];
            n_Body_y[2999] = c_Body_y[2999];
            n_Body_x[3000] = c_Body_x[3000];
            n_Body_y[3000] = c_Body_y[3000];
            n_Body_x[3001] = c_Body_x[3001];
            n_Body_y[3001] = c_Body_y[3001];
            n_Body_x[3002] = c_Body_x[3002];
            n_Body_y[3002] = c_Body_y[3002];
            n_Body_x[3003] = c_Body_x[3003];
            n_Body_y[3003] = c_Body_y[3003];
            n_Body_x[3004] = c_Body_x[3004];
            n_Body_y[3004] = c_Body_y[3004];
            n_Body_x[3005] = c_Body_x[3005];
            n_Body_y[3005] = c_Body_y[3005];
            n_Body_x[3006] = c_Body_x[3006];
            n_Body_y[3006] = c_Body_y[3006];
            n_Body_x[3007] = c_Body_x[3007];
            n_Body_y[3007] = c_Body_y[3007];
            n_Body_x[3008] = c_Body_x[3008];
            n_Body_y[3008] = c_Body_y[3008];
            n_Body_x[3009] = c_Body_x[3009];
            n_Body_y[3009] = c_Body_y[3009];
            n_Body_x[3010] = c_Body_x[3010];
            n_Body_y[3010] = c_Body_y[3010];
            n_Body_x[3011] = c_Body_x[3011];
            n_Body_y[3011] = c_Body_y[3011];
            n_Body_x[3012] = c_Body_x[3012];
            n_Body_y[3012] = c_Body_y[3012];
            n_Body_x[3013] = c_Body_x[3013];
            n_Body_y[3013] = c_Body_y[3013];
            n_Body_x[3014] = c_Body_x[3014];
            n_Body_y[3014] = c_Body_y[3014];
            n_Body_x[3015] = c_Body_x[3015];
            n_Body_y[3015] = c_Body_y[3015];
            n_Body_x[3016] = c_Body_x[3016];
            n_Body_y[3016] = c_Body_y[3016];
            n_Body_x[3017] = c_Body_x[3017];
            n_Body_y[3017] = c_Body_y[3017];
            n_Body_x[3018] = c_Body_x[3018];
            n_Body_y[3018] = c_Body_y[3018];
            n_Body_x[3019] = c_Body_x[3019];
            n_Body_y[3019] = c_Body_y[3019];
            n_Body_x[3020] = c_Body_x[3020];
            n_Body_y[3020] = c_Body_y[3020];
            n_Body_x[3021] = c_Body_x[3021];
            n_Body_y[3021] = c_Body_y[3021];
            n_Body_x[3022] = c_Body_x[3022];
            n_Body_y[3022] = c_Body_y[3022];
            n_Body_x[3023] = c_Body_x[3023];
            n_Body_y[3023] = c_Body_y[3023];
            n_Body_x[3024] = c_Body_x[3024];
            n_Body_y[3024] = c_Body_y[3024];
            n_Body_x[3025] = c_Body_x[3025];
            n_Body_y[3025] = c_Body_y[3025];
            n_Body_x[3026] = c_Body_x[3026];
            n_Body_y[3026] = c_Body_y[3026];
            n_Body_x[3027] = c_Body_x[3027];
            n_Body_y[3027] = c_Body_y[3027];
            n_Body_x[3028] = c_Body_x[3028];
            n_Body_y[3028] = c_Body_y[3028];
            n_Body_x[3029] = c_Body_x[3029];
            n_Body_y[3029] = c_Body_y[3029];
            n_Body_x[3030] = c_Body_x[3030];
            n_Body_y[3030] = c_Body_y[3030];
            n_Body_x[3031] = c_Body_x[3031];
            n_Body_y[3031] = c_Body_y[3031];
            n_Body_x[3032] = c_Body_x[3032];
            n_Body_y[3032] = c_Body_y[3032];
            n_Body_x[3033] = c_Body_x[3033];
            n_Body_y[3033] = c_Body_y[3033];
            n_Body_x[3034] = c_Body_x[3034];
            n_Body_y[3034] = c_Body_y[3034];
            n_Body_x[3035] = c_Body_x[3035];
            n_Body_y[3035] = c_Body_y[3035];
            n_Body_x[3036] = c_Body_x[3036];
            n_Body_y[3036] = c_Body_y[3036];
            n_Body_x[3037] = c_Body_x[3037];
            n_Body_y[3037] = c_Body_y[3037];
            n_Body_x[3038] = c_Body_x[3038];
            n_Body_y[3038] = c_Body_y[3038];
            n_Body_x[3039] = c_Body_x[3039];
            n_Body_y[3039] = c_Body_y[3039];
            n_Body_x[3040] = c_Body_x[3040];
            n_Body_y[3040] = c_Body_y[3040];
            n_Body_x[3041] = c_Body_x[3041];
            n_Body_y[3041] = c_Body_y[3041];
            n_Body_x[3042] = c_Body_x[3042];
            n_Body_y[3042] = c_Body_y[3042];
            n_Body_x[3043] = c_Body_x[3043];
            n_Body_y[3043] = c_Body_y[3043];
            n_Body_x[3044] = c_Body_x[3044];
            n_Body_y[3044] = c_Body_y[3044];
            n_Body_x[3045] = c_Body_x[3045];
            n_Body_y[3045] = c_Body_y[3045];
            n_Body_x[3046] = c_Body_x[3046];
            n_Body_y[3046] = c_Body_y[3046];
            n_Body_x[3047] = c_Body_x[3047];
            n_Body_y[3047] = c_Body_y[3047];
            n_Body_x[3048] = c_Body_x[3048];
            n_Body_y[3048] = c_Body_y[3048];
            n_Body_x[3049] = c_Body_x[3049];
            n_Body_y[3049] = c_Body_y[3049];
            n_Body_x[3050] = c_Body_x[3050];
            n_Body_y[3050] = c_Body_y[3050];
            n_Body_x[3051] = c_Body_x[3051];
            n_Body_y[3051] = c_Body_y[3051];
            n_Body_x[3052] = c_Body_x[3052];
            n_Body_y[3052] = c_Body_y[3052];
            n_Body_x[3053] = c_Body_x[3053];
            n_Body_y[3053] = c_Body_y[3053];
            n_Body_x[3054] = c_Body_x[3054];
            n_Body_y[3054] = c_Body_y[3054];
            n_Body_x[3055] = c_Body_x[3055];
            n_Body_y[3055] = c_Body_y[3055];
            n_Body_x[3056] = c_Body_x[3056];
            n_Body_y[3056] = c_Body_y[3056];
            n_Body_x[3057] = c_Body_x[3057];
            n_Body_y[3057] = c_Body_y[3057];
            n_Body_x[3058] = c_Body_x[3058];
            n_Body_y[3058] = c_Body_y[3058];
            n_Body_x[3059] = c_Body_x[3059];
            n_Body_y[3059] = c_Body_y[3059];
            n_Body_x[3060] = c_Body_x[3060];
            n_Body_y[3060] = c_Body_y[3060];
            n_Body_x[3061] = c_Body_x[3061];
            n_Body_y[3061] = c_Body_y[3061];
            n_Body_x[3062] = c_Body_x[3062];
            n_Body_y[3062] = c_Body_y[3062];
            n_Body_x[3063] = c_Body_x[3063];
            n_Body_y[3063] = c_Body_y[3063];
            n_Body_x[3064] = c_Body_x[3064];
            n_Body_y[3064] = c_Body_y[3064];
            n_Body_x[3065] = c_Body_x[3065];
            n_Body_y[3065] = c_Body_y[3065];
            n_Body_x[3066] = c_Body_x[3066];
            n_Body_y[3066] = c_Body_y[3066];
            n_Body_x[3067] = c_Body_x[3067];
            n_Body_y[3067] = c_Body_y[3067];
            n_Body_x[3068] = c_Body_x[3068];
            n_Body_y[3068] = c_Body_y[3068];
            n_Body_x[3069] = c_Body_x[3069];
            n_Body_y[3069] = c_Body_y[3069];
            n_Body_x[3070] = c_Body_x[3070];
            n_Body_y[3070] = c_Body_y[3070];
            n_Body_x[3071] = c_Body_x[3071];
            n_Body_y[3071] = c_Body_y[3071];

        case(c_State)
            IDLE : begin
                n_ClkCnt = c_ClkCnt + 1;
                if(!(&i_Push)) begin
                    n_State = RUN;
                    n_ClkCnt = 0;
                end
            end
            RUN  : begin
                n_ClkCnt = isLstClk ? 0 : c_ClkCnt + c_Speed;
                n_Push = !i_Push[0] ? 0 :
                         !i_Push[1] ? 1 :
                         !i_Push[2] ? 2 :
                         !i_Push[3] ? 3 : c_Push;

                if(isLstClk) begin
                    //속도 조절 로직
                    n_SpdTimeCnt = isSpdDw ? 0 : c_SpdTimeCnt + 1;
                    n_Speed = isSpdDw ? DEF_SPD : c_Speed; // 시간 다되면 기본 속도

                    //헤드 위치, 방향 갱신
                    {n_Head_x,n_Head_y} = {SH_o_Head_x,SH_o_Head_y};
                    n_Way = SH_o_Way;

                    n_State = CHANGE;
                end
                n_State = i_Pause ? PAUSE : RUN;
            end
            CHANGE : begin // n_Head값들 바뀐거로 사이즈값 변경이랑 게임 오버 판정, 아이템 새로 만듬
                if(isEat) begin
                    n_Size = c_Size + (c_Speed >> 1); // 속도의 절반만큼 점수가 오름
                    //n_Item_x = ;
                    //n_Item_y = ; 
                    n_Speed = c_Speed + 1;
                    n_SpdTimeCnt = 0;
                end
                n_State = o_isMakeItem_Done ? (isGameOver ? STOP : SETBODY) : c_State;
            end
            SETBODY : begin // 사이즈값 갱신했으니 그걸로 몸통 큐 갱신
                n_Body_x[0] = c_Head_x;
                n_Body_y[0] = c_Head_y;
                
                //무수히 많은 if-else문들...
                    if (n_Size > 1) begin
                        n_Body_x[1] = c_Body_x[0];
                        n_Body_y[1] = c_Body_y[0];
                    end else begin
                        n_Body_x[1] = c_Body_x[c_Size-1];
                        n_Body_y[1] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2) begin
                        n_Body_x[2] = c_Body_x[1];
                        n_Body_y[2] = c_Body_y[1];
                    end else begin
                        n_Body_x[2] = c_Body_x[c_Size-1];
                        n_Body_y[2] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3) begin
                        n_Body_x[3] = c_Body_x[2];
                        n_Body_y[3] = c_Body_y[2];
                    end else begin
                        n_Body_x[3] = c_Body_x[c_Size-1];
                        n_Body_y[3] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 4) begin
                        n_Body_x[4] = c_Body_x[3];
                        n_Body_y[4] = c_Body_y[3];
                    end else begin
                        n_Body_x[4] = c_Body_x[c_Size-1];
                        n_Body_y[4] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 5) begin
                        n_Body_x[5] = c_Body_x[4];
                        n_Body_y[5] = c_Body_y[4];
                    end else begin
                        n_Body_x[5] = c_Body_x[c_Size-1];
                        n_Body_y[5] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 6) begin
                        n_Body_x[6] = c_Body_x[5];
                        n_Body_y[6] = c_Body_y[5];
                    end else begin
                        n_Body_x[6] = c_Body_x[c_Size-1];
                        n_Body_y[6] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 7) begin
                        n_Body_x[7] = c_Body_x[6];
                        n_Body_y[7] = c_Body_y[6];
                    end else begin
                        n_Body_x[7] = c_Body_x[c_Size-1];
                        n_Body_y[7] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 8) begin
                        n_Body_x[8] = c_Body_x[7];
                        n_Body_y[8] = c_Body_y[7];
                    end else begin
                        n_Body_x[8] = c_Body_x[c_Size-1];
                        n_Body_y[8] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 9) begin
                        n_Body_x[9] = c_Body_x[8];
                        n_Body_y[9] = c_Body_y[8];
                    end else begin
                        n_Body_x[9] = c_Body_x[c_Size-1];
                        n_Body_y[9] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 10) begin
                        n_Body_x[10] = c_Body_x[9];
                        n_Body_y[10] = c_Body_y[9];
                    end else begin
                        n_Body_x[10] = c_Body_x[c_Size-1];
                        n_Body_y[10] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 11) begin
                        n_Body_x[11] = c_Body_x[10];
                        n_Body_y[11] = c_Body_y[10];
                    end else begin
                        n_Body_x[11] = c_Body_x[c_Size-1];
                        n_Body_y[11] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 12) begin
                        n_Body_x[12] = c_Body_x[11];
                        n_Body_y[12] = c_Body_y[11];
                    end else begin
                        n_Body_x[12] = c_Body_x[c_Size-1];
                        n_Body_y[12] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 13) begin
                        n_Body_x[13] = c_Body_x[12];
                        n_Body_y[13] = c_Body_y[12];
                    end else begin
                        n_Body_x[13] = c_Body_x[c_Size-1];
                        n_Body_y[13] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 14) begin
                        n_Body_x[14] = c_Body_x[13];
                        n_Body_y[14] = c_Body_y[13];
                    end else begin
                        n_Body_x[14] = c_Body_x[c_Size-1];
                        n_Body_y[14] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 15) begin
                        n_Body_x[15] = c_Body_x[14];
                        n_Body_y[15] = c_Body_y[14];
                    end else begin
                        n_Body_x[15] = c_Body_x[c_Size-1];
                        n_Body_y[15] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 16) begin
                        n_Body_x[16] = c_Body_x[15];
                        n_Body_y[16] = c_Body_y[15];
                    end else begin
                        n_Body_x[16] = c_Body_x[c_Size-1];
                        n_Body_y[16] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 17) begin
                        n_Body_x[17] = c_Body_x[16];
                        n_Body_y[17] = c_Body_y[16];
                    end else begin
                        n_Body_x[17] = c_Body_x[c_Size-1];
                        n_Body_y[17] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 18) begin
                        n_Body_x[18] = c_Body_x[17];
                        n_Body_y[18] = c_Body_y[17];
                    end else begin
                        n_Body_x[18] = c_Body_x[c_Size-1];
                        n_Body_y[18] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 19) begin
                        n_Body_x[19] = c_Body_x[18];
                        n_Body_y[19] = c_Body_y[18];
                    end else begin
                        n_Body_x[19] = c_Body_x[c_Size-1];
                        n_Body_y[19] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 20) begin
                        n_Body_x[20] = c_Body_x[19];
                        n_Body_y[20] = c_Body_y[19];
                    end else begin
                        n_Body_x[20] = c_Body_x[c_Size-1];
                        n_Body_y[20] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 21) begin
                        n_Body_x[21] = c_Body_x[20];
                        n_Body_y[21] = c_Body_y[20];
                    end else begin
                        n_Body_x[21] = c_Body_x[c_Size-1];
                        n_Body_y[21] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 22) begin
                        n_Body_x[22] = c_Body_x[21];
                        n_Body_y[22] = c_Body_y[21];
                    end else begin
                        n_Body_x[22] = c_Body_x[c_Size-1];
                        n_Body_y[22] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 23) begin
                        n_Body_x[23] = c_Body_x[22];
                        n_Body_y[23] = c_Body_y[22];
                    end else begin
                        n_Body_x[23] = c_Body_x[c_Size-1];
                        n_Body_y[23] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 24) begin
                        n_Body_x[24] = c_Body_x[23];
                        n_Body_y[24] = c_Body_y[23];
                    end else begin
                        n_Body_x[24] = c_Body_x[c_Size-1];
                        n_Body_y[24] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 25) begin
                        n_Body_x[25] = c_Body_x[24];
                        n_Body_y[25] = c_Body_y[24];
                    end else begin
                        n_Body_x[25] = c_Body_x[c_Size-1];
                        n_Body_y[25] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 26) begin
                        n_Body_x[26] = c_Body_x[25];
                        n_Body_y[26] = c_Body_y[25];
                    end else begin
                        n_Body_x[26] = c_Body_x[c_Size-1];
                        n_Body_y[26] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 27) begin
                        n_Body_x[27] = c_Body_x[26];
                        n_Body_y[27] = c_Body_y[26];
                    end else begin
                        n_Body_x[27] = c_Body_x[c_Size-1];
                        n_Body_y[27] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 28) begin
                        n_Body_x[28] = c_Body_x[27];
                        n_Body_y[28] = c_Body_y[27];
                    end else begin
                        n_Body_x[28] = c_Body_x[c_Size-1];
                        n_Body_y[28] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 29) begin
                        n_Body_x[29] = c_Body_x[28];
                        n_Body_y[29] = c_Body_y[28];
                    end else begin
                        n_Body_x[29] = c_Body_x[c_Size-1];
                        n_Body_y[29] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 30) begin
                        n_Body_x[30] = c_Body_x[29];
                        n_Body_y[30] = c_Body_y[29];
                    end else begin
                        n_Body_x[30] = c_Body_x[c_Size-1];
                        n_Body_y[30] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 31) begin
                        n_Body_x[31] = c_Body_x[30];
                        n_Body_y[31] = c_Body_y[30];
                    end else begin
                        n_Body_x[31] = c_Body_x[c_Size-1];
                        n_Body_y[31] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 32) begin
                        n_Body_x[32] = c_Body_x[31];
                        n_Body_y[32] = c_Body_y[31];
                    end else begin
                        n_Body_x[32] = c_Body_x[c_Size-1];
                        n_Body_y[32] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 33) begin
                        n_Body_x[33] = c_Body_x[32];
                        n_Body_y[33] = c_Body_y[32];
                    end else begin
                        n_Body_x[33] = c_Body_x[c_Size-1];
                        n_Body_y[33] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 34) begin
                        n_Body_x[34] = c_Body_x[33];
                        n_Body_y[34] = c_Body_y[33];
                    end else begin
                        n_Body_x[34] = c_Body_x[c_Size-1];
                        n_Body_y[34] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 35) begin
                        n_Body_x[35] = c_Body_x[34];
                        n_Body_y[35] = c_Body_y[34];
                    end else begin
                        n_Body_x[35] = c_Body_x[c_Size-1];
                        n_Body_y[35] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 36) begin
                        n_Body_x[36] = c_Body_x[35];
                        n_Body_y[36] = c_Body_y[35];
                    end else begin
                        n_Body_x[36] = c_Body_x[c_Size-1];
                        n_Body_y[36] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 37) begin
                        n_Body_x[37] = c_Body_x[36];
                        n_Body_y[37] = c_Body_y[36];
                    end else begin
                        n_Body_x[37] = c_Body_x[c_Size-1];
                        n_Body_y[37] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 38) begin
                        n_Body_x[38] = c_Body_x[37];
                        n_Body_y[38] = c_Body_y[37];
                    end else begin
                        n_Body_x[38] = c_Body_x[c_Size-1];
                        n_Body_y[38] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 39) begin
                        n_Body_x[39] = c_Body_x[38];
                        n_Body_y[39] = c_Body_y[38];
                    end else begin
                        n_Body_x[39] = c_Body_x[c_Size-1];
                        n_Body_y[39] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 40) begin
                        n_Body_x[40] = c_Body_x[39];
                        n_Body_y[40] = c_Body_y[39];
                    end else begin
                        n_Body_x[40] = c_Body_x[c_Size-1];
                        n_Body_y[40] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 41) begin
                        n_Body_x[41] = c_Body_x[40];
                        n_Body_y[41] = c_Body_y[40];
                    end else begin
                        n_Body_x[41] = c_Body_x[c_Size-1];
                        n_Body_y[41] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 42) begin
                        n_Body_x[42] = c_Body_x[41];
                        n_Body_y[42] = c_Body_y[41];
                    end else begin
                        n_Body_x[42] = c_Body_x[c_Size-1];
                        n_Body_y[42] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 43) begin
                        n_Body_x[43] = c_Body_x[42];
                        n_Body_y[43] = c_Body_y[42];
                    end else begin
                        n_Body_x[43] = c_Body_x[c_Size-1];
                        n_Body_y[43] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 44) begin
                        n_Body_x[44] = c_Body_x[43];
                        n_Body_y[44] = c_Body_y[43];
                    end else begin
                        n_Body_x[44] = c_Body_x[c_Size-1];
                        n_Body_y[44] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 45) begin
                        n_Body_x[45] = c_Body_x[44];
                        n_Body_y[45] = c_Body_y[44];
                    end else begin
                        n_Body_x[45] = c_Body_x[c_Size-1];
                        n_Body_y[45] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 46) begin
                        n_Body_x[46] = c_Body_x[45];
                        n_Body_y[46] = c_Body_y[45];
                    end else begin
                        n_Body_x[46] = c_Body_x[c_Size-1];
                        n_Body_y[46] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 47) begin
                        n_Body_x[47] = c_Body_x[46];
                        n_Body_y[47] = c_Body_y[46];
                    end else begin
                        n_Body_x[47] = c_Body_x[c_Size-1];
                        n_Body_y[47] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 48) begin
                        n_Body_x[48] = c_Body_x[47];
                        n_Body_y[48] = c_Body_y[47];
                    end else begin
                        n_Body_x[48] = c_Body_x[c_Size-1];
                        n_Body_y[48] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 49) begin
                        n_Body_x[49] = c_Body_x[48];
                        n_Body_y[49] = c_Body_y[48];
                    end else begin
                        n_Body_x[49] = c_Body_x[c_Size-1];
                        n_Body_y[49] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 50) begin
                        n_Body_x[50] = c_Body_x[49];
                        n_Body_y[50] = c_Body_y[49];
                    end else begin
                        n_Body_x[50] = c_Body_x[c_Size-1];
                        n_Body_y[50] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 51) begin
                        n_Body_x[51] = c_Body_x[50];
                        n_Body_y[51] = c_Body_y[50];
                    end else begin
                        n_Body_x[51] = c_Body_x[c_Size-1];
                        n_Body_y[51] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 52) begin
                        n_Body_x[52] = c_Body_x[51];
                        n_Body_y[52] = c_Body_y[51];
                    end else begin
                        n_Body_x[52] = c_Body_x[c_Size-1];
                        n_Body_y[52] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 53) begin
                        n_Body_x[53] = c_Body_x[52];
                        n_Body_y[53] = c_Body_y[52];
                    end else begin
                        n_Body_x[53] = c_Body_x[c_Size-1];
                        n_Body_y[53] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 54) begin
                        n_Body_x[54] = c_Body_x[53];
                        n_Body_y[54] = c_Body_y[53];
                    end else begin
                        n_Body_x[54] = c_Body_x[c_Size-1];
                        n_Body_y[54] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 55) begin
                        n_Body_x[55] = c_Body_x[54];
                        n_Body_y[55] = c_Body_y[54];
                    end else begin
                        n_Body_x[55] = c_Body_x[c_Size-1];
                        n_Body_y[55] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 56) begin
                        n_Body_x[56] = c_Body_x[55];
                        n_Body_y[56] = c_Body_y[55];
                    end else begin
                        n_Body_x[56] = c_Body_x[c_Size-1];
                        n_Body_y[56] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 57) begin
                        n_Body_x[57] = c_Body_x[56];
                        n_Body_y[57] = c_Body_y[56];
                    end else begin
                        n_Body_x[57] = c_Body_x[c_Size-1];
                        n_Body_y[57] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 58) begin
                        n_Body_x[58] = c_Body_x[57];
                        n_Body_y[58] = c_Body_y[57];
                    end else begin
                        n_Body_x[58] = c_Body_x[c_Size-1];
                        n_Body_y[58] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 59) begin
                        n_Body_x[59] = c_Body_x[58];
                        n_Body_y[59] = c_Body_y[58];
                    end else begin
                        n_Body_x[59] = c_Body_x[c_Size-1];
                        n_Body_y[59] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 60) begin
                        n_Body_x[60] = c_Body_x[59];
                        n_Body_y[60] = c_Body_y[59];
                    end else begin
                        n_Body_x[60] = c_Body_x[c_Size-1];
                        n_Body_y[60] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 61) begin
                        n_Body_x[61] = c_Body_x[60];
                        n_Body_y[61] = c_Body_y[60];
                    end else begin
                        n_Body_x[61] = c_Body_x[c_Size-1];
                        n_Body_y[61] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 62) begin
                        n_Body_x[62] = c_Body_x[61];
                        n_Body_y[62] = c_Body_y[61];
                    end else begin
                        n_Body_x[62] = c_Body_x[c_Size-1];
                        n_Body_y[62] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 63) begin
                        n_Body_x[63] = c_Body_x[62];
                        n_Body_y[63] = c_Body_y[62];
                    end else begin
                        n_Body_x[63] = c_Body_x[c_Size-1];
                        n_Body_y[63] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 64) begin
                        n_Body_x[64] = c_Body_x[63];
                        n_Body_y[64] = c_Body_y[63];
                    end else begin
                        n_Body_x[64] = c_Body_x[c_Size-1];
                        n_Body_y[64] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 65) begin
                        n_Body_x[65] = c_Body_x[64];
                        n_Body_y[65] = c_Body_y[64];
                    end else begin
                        n_Body_x[65] = c_Body_x[c_Size-1];
                        n_Body_y[65] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 66) begin
                        n_Body_x[66] = c_Body_x[65];
                        n_Body_y[66] = c_Body_y[65];
                    end else begin
                        n_Body_x[66] = c_Body_x[c_Size-1];
                        n_Body_y[66] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 67) begin
                        n_Body_x[67] = c_Body_x[66];
                        n_Body_y[67] = c_Body_y[66];
                    end else begin
                        n_Body_x[67] = c_Body_x[c_Size-1];
                        n_Body_y[67] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 68) begin
                        n_Body_x[68] = c_Body_x[67];
                        n_Body_y[68] = c_Body_y[67];
                    end else begin
                        n_Body_x[68] = c_Body_x[c_Size-1];
                        n_Body_y[68] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 69) begin
                        n_Body_x[69] = c_Body_x[68];
                        n_Body_y[69] = c_Body_y[68];
                    end else begin
                        n_Body_x[69] = c_Body_x[c_Size-1];
                        n_Body_y[69] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 70) begin
                        n_Body_x[70] = c_Body_x[69];
                        n_Body_y[70] = c_Body_y[69];
                    end else begin
                        n_Body_x[70] = c_Body_x[c_Size-1];
                        n_Body_y[70] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 71) begin
                        n_Body_x[71] = c_Body_x[70];
                        n_Body_y[71] = c_Body_y[70];
                    end else begin
                        n_Body_x[71] = c_Body_x[c_Size-1];
                        n_Body_y[71] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 72) begin
                        n_Body_x[72] = c_Body_x[71];
                        n_Body_y[72] = c_Body_y[71];
                    end else begin
                        n_Body_x[72] = c_Body_x[c_Size-1];
                        n_Body_y[72] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 73) begin
                        n_Body_x[73] = c_Body_x[72];
                        n_Body_y[73] = c_Body_y[72];
                    end else begin
                        n_Body_x[73] = c_Body_x[c_Size-1];
                        n_Body_y[73] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 74) begin
                        n_Body_x[74] = c_Body_x[73];
                        n_Body_y[74] = c_Body_y[73];
                    end else begin
                        n_Body_x[74] = c_Body_x[c_Size-1];
                        n_Body_y[74] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 75) begin
                        n_Body_x[75] = c_Body_x[74];
                        n_Body_y[75] = c_Body_y[74];
                    end else begin
                        n_Body_x[75] = c_Body_x[c_Size-1];
                        n_Body_y[75] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 76) begin
                        n_Body_x[76] = c_Body_x[75];
                        n_Body_y[76] = c_Body_y[75];
                    end else begin
                        n_Body_x[76] = c_Body_x[c_Size-1];
                        n_Body_y[76] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 77) begin
                        n_Body_x[77] = c_Body_x[76];
                        n_Body_y[77] = c_Body_y[76];
                    end else begin
                        n_Body_x[77] = c_Body_x[c_Size-1];
                        n_Body_y[77] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 78) begin
                        n_Body_x[78] = c_Body_x[77];
                        n_Body_y[78] = c_Body_y[77];
                    end else begin
                        n_Body_x[78] = c_Body_x[c_Size-1];
                        n_Body_y[78] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 79) begin
                        n_Body_x[79] = c_Body_x[78];
                        n_Body_y[79] = c_Body_y[78];
                    end else begin
                        n_Body_x[79] = c_Body_x[c_Size-1];
                        n_Body_y[79] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 80) begin
                        n_Body_x[80] = c_Body_x[79];
                        n_Body_y[80] = c_Body_y[79];
                    end else begin
                        n_Body_x[80] = c_Body_x[c_Size-1];
                        n_Body_y[80] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 81) begin
                        n_Body_x[81] = c_Body_x[80];
                        n_Body_y[81] = c_Body_y[80];
                    end else begin
                        n_Body_x[81] = c_Body_x[c_Size-1];
                        n_Body_y[81] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 82) begin
                        n_Body_x[82] = c_Body_x[81];
                        n_Body_y[82] = c_Body_y[81];
                    end else begin
                        n_Body_x[82] = c_Body_x[c_Size-1];
                        n_Body_y[82] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 83) begin
                        n_Body_x[83] = c_Body_x[82];
                        n_Body_y[83] = c_Body_y[82];
                    end else begin
                        n_Body_x[83] = c_Body_x[c_Size-1];
                        n_Body_y[83] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 84) begin
                        n_Body_x[84] = c_Body_x[83];
                        n_Body_y[84] = c_Body_y[83];
                    end else begin
                        n_Body_x[84] = c_Body_x[c_Size-1];
                        n_Body_y[84] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 85) begin
                        n_Body_x[85] = c_Body_x[84];
                        n_Body_y[85] = c_Body_y[84];
                    end else begin
                        n_Body_x[85] = c_Body_x[c_Size-1];
                        n_Body_y[85] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 86) begin
                        n_Body_x[86] = c_Body_x[85];
                        n_Body_y[86] = c_Body_y[85];
                    end else begin
                        n_Body_x[86] = c_Body_x[c_Size-1];
                        n_Body_y[86] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 87) begin
                        n_Body_x[87] = c_Body_x[86];
                        n_Body_y[87] = c_Body_y[86];
                    end else begin
                        n_Body_x[87] = c_Body_x[c_Size-1];
                        n_Body_y[87] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 88) begin
                        n_Body_x[88] = c_Body_x[87];
                        n_Body_y[88] = c_Body_y[87];
                    end else begin
                        n_Body_x[88] = c_Body_x[c_Size-1];
                        n_Body_y[88] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 89) begin
                        n_Body_x[89] = c_Body_x[88];
                        n_Body_y[89] = c_Body_y[88];
                    end else begin
                        n_Body_x[89] = c_Body_x[c_Size-1];
                        n_Body_y[89] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 90) begin
                        n_Body_x[90] = c_Body_x[89];
                        n_Body_y[90] = c_Body_y[89];
                    end else begin
                        n_Body_x[90] = c_Body_x[c_Size-1];
                        n_Body_y[90] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 91) begin
                        n_Body_x[91] = c_Body_x[90];
                        n_Body_y[91] = c_Body_y[90];
                    end else begin
                        n_Body_x[91] = c_Body_x[c_Size-1];
                        n_Body_y[91] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 92) begin
                        n_Body_x[92] = c_Body_x[91];
                        n_Body_y[92] = c_Body_y[91];
                    end else begin
                        n_Body_x[92] = c_Body_x[c_Size-1];
                        n_Body_y[92] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 93) begin
                        n_Body_x[93] = c_Body_x[92];
                        n_Body_y[93] = c_Body_y[92];
                    end else begin
                        n_Body_x[93] = c_Body_x[c_Size-1];
                        n_Body_y[93] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 94) begin
                        n_Body_x[94] = c_Body_x[93];
                        n_Body_y[94] = c_Body_y[93];
                    end else begin
                        n_Body_x[94] = c_Body_x[c_Size-1];
                        n_Body_y[94] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 95) begin
                        n_Body_x[95] = c_Body_x[94];
                        n_Body_y[95] = c_Body_y[94];
                    end else begin
                        n_Body_x[95] = c_Body_x[c_Size-1];
                        n_Body_y[95] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 96) begin
                        n_Body_x[96] = c_Body_x[95];
                        n_Body_y[96] = c_Body_y[95];
                    end else begin
                        n_Body_x[96] = c_Body_x[c_Size-1];
                        n_Body_y[96] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 97) begin
                        n_Body_x[97] = c_Body_x[96];
                        n_Body_y[97] = c_Body_y[96];
                    end else begin
                        n_Body_x[97] = c_Body_x[c_Size-1];
                        n_Body_y[97] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 98) begin
                        n_Body_x[98] = c_Body_x[97];
                        n_Body_y[98] = c_Body_y[97];
                    end else begin
                        n_Body_x[98] = c_Body_x[c_Size-1];
                        n_Body_y[98] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 99) begin
                        n_Body_x[99] = c_Body_x[98];
                        n_Body_y[99] = c_Body_y[98];
                    end else begin
                        n_Body_x[99] = c_Body_x[c_Size-1];
                        n_Body_y[99] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 100) begin
                        n_Body_x[100] = c_Body_x[99];
                        n_Body_y[100] = c_Body_y[99];
                    end else begin
                        n_Body_x[100] = c_Body_x[c_Size-1];
                        n_Body_y[100] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 101) begin
                        n_Body_x[101] = c_Body_x[100];
                        n_Body_y[101] = c_Body_y[100];
                    end else begin
                        n_Body_x[101] = c_Body_x[c_Size-1];
                        n_Body_y[101] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 102) begin
                        n_Body_x[102] = c_Body_x[101];
                        n_Body_y[102] = c_Body_y[101];
                    end else begin
                        n_Body_x[102] = c_Body_x[c_Size-1];
                        n_Body_y[102] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 103) begin
                        n_Body_x[103] = c_Body_x[102];
                        n_Body_y[103] = c_Body_y[102];
                    end else begin
                        n_Body_x[103] = c_Body_x[c_Size-1];
                        n_Body_y[103] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 104) begin
                        n_Body_x[104] = c_Body_x[103];
                        n_Body_y[104] = c_Body_y[103];
                    end else begin
                        n_Body_x[104] = c_Body_x[c_Size-1];
                        n_Body_y[104] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 105) begin
                        n_Body_x[105] = c_Body_x[104];
                        n_Body_y[105] = c_Body_y[104];
                    end else begin
                        n_Body_x[105] = c_Body_x[c_Size-1];
                        n_Body_y[105] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 106) begin
                        n_Body_x[106] = c_Body_x[105];
                        n_Body_y[106] = c_Body_y[105];
                    end else begin
                        n_Body_x[106] = c_Body_x[c_Size-1];
                        n_Body_y[106] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 107) begin
                        n_Body_x[107] = c_Body_x[106];
                        n_Body_y[107] = c_Body_y[106];
                    end else begin
                        n_Body_x[107] = c_Body_x[c_Size-1];
                        n_Body_y[107] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 108) begin
                        n_Body_x[108] = c_Body_x[107];
                        n_Body_y[108] = c_Body_y[107];
                    end else begin
                        n_Body_x[108] = c_Body_x[c_Size-1];
                        n_Body_y[108] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 109) begin
                        n_Body_x[109] = c_Body_x[108];
                        n_Body_y[109] = c_Body_y[108];
                    end else begin
                        n_Body_x[109] = c_Body_x[c_Size-1];
                        n_Body_y[109] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 110) begin
                        n_Body_x[110] = c_Body_x[109];
                        n_Body_y[110] = c_Body_y[109];
                    end else begin
                        n_Body_x[110] = c_Body_x[c_Size-1];
                        n_Body_y[110] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 111) begin
                        n_Body_x[111] = c_Body_x[110];
                        n_Body_y[111] = c_Body_y[110];
                    end else begin
                        n_Body_x[111] = c_Body_x[c_Size-1];
                        n_Body_y[111] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 112) begin
                        n_Body_x[112] = c_Body_x[111];
                        n_Body_y[112] = c_Body_y[111];
                    end else begin
                        n_Body_x[112] = c_Body_x[c_Size-1];
                        n_Body_y[112] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 113) begin
                        n_Body_x[113] = c_Body_x[112];
                        n_Body_y[113] = c_Body_y[112];
                    end else begin
                        n_Body_x[113] = c_Body_x[c_Size-1];
                        n_Body_y[113] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 114) begin
                        n_Body_x[114] = c_Body_x[113];
                        n_Body_y[114] = c_Body_y[113];
                    end else begin
                        n_Body_x[114] = c_Body_x[c_Size-1];
                        n_Body_y[114] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 115) begin
                        n_Body_x[115] = c_Body_x[114];
                        n_Body_y[115] = c_Body_y[114];
                    end else begin
                        n_Body_x[115] = c_Body_x[c_Size-1];
                        n_Body_y[115] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 116) begin
                        n_Body_x[116] = c_Body_x[115];
                        n_Body_y[116] = c_Body_y[115];
                    end else begin
                        n_Body_x[116] = c_Body_x[c_Size-1];
                        n_Body_y[116] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 117) begin
                        n_Body_x[117] = c_Body_x[116];
                        n_Body_y[117] = c_Body_y[116];
                    end else begin
                        n_Body_x[117] = c_Body_x[c_Size-1];
                        n_Body_y[117] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 118) begin
                        n_Body_x[118] = c_Body_x[117];
                        n_Body_y[118] = c_Body_y[117];
                    end else begin
                        n_Body_x[118] = c_Body_x[c_Size-1];
                        n_Body_y[118] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 119) begin
                        n_Body_x[119] = c_Body_x[118];
                        n_Body_y[119] = c_Body_y[118];
                    end else begin
                        n_Body_x[119] = c_Body_x[c_Size-1];
                        n_Body_y[119] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 120) begin
                        n_Body_x[120] = c_Body_x[119];
                        n_Body_y[120] = c_Body_y[119];
                    end else begin
                        n_Body_x[120] = c_Body_x[c_Size-1];
                        n_Body_y[120] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 121) begin
                        n_Body_x[121] = c_Body_x[120];
                        n_Body_y[121] = c_Body_y[120];
                    end else begin
                        n_Body_x[121] = c_Body_x[c_Size-1];
                        n_Body_y[121] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 122) begin
                        n_Body_x[122] = c_Body_x[121];
                        n_Body_y[122] = c_Body_y[121];
                    end else begin
                        n_Body_x[122] = c_Body_x[c_Size-1];
                        n_Body_y[122] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 123) begin
                        n_Body_x[123] = c_Body_x[122];
                        n_Body_y[123] = c_Body_y[122];
                    end else begin
                        n_Body_x[123] = c_Body_x[c_Size-1];
                        n_Body_y[123] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 124) begin
                        n_Body_x[124] = c_Body_x[123];
                        n_Body_y[124] = c_Body_y[123];
                    end else begin
                        n_Body_x[124] = c_Body_x[c_Size-1];
                        n_Body_y[124] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 125) begin
                        n_Body_x[125] = c_Body_x[124];
                        n_Body_y[125] = c_Body_y[124];
                    end else begin
                        n_Body_x[125] = c_Body_x[c_Size-1];
                        n_Body_y[125] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 126) begin
                        n_Body_x[126] = c_Body_x[125];
                        n_Body_y[126] = c_Body_y[125];
                    end else begin
                        n_Body_x[126] = c_Body_x[c_Size-1];
                        n_Body_y[126] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 127) begin
                        n_Body_x[127] = c_Body_x[126];
                        n_Body_y[127] = c_Body_y[126];
                    end else begin
                        n_Body_x[127] = c_Body_x[c_Size-1];
                        n_Body_y[127] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 128) begin
                        n_Body_x[128] = c_Body_x[127];
                        n_Body_y[128] = c_Body_y[127];
                    end else begin
                        n_Body_x[128] = c_Body_x[c_Size-1];
                        n_Body_y[128] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 129) begin
                        n_Body_x[129] = c_Body_x[128];
                        n_Body_y[129] = c_Body_y[128];
                    end else begin
                        n_Body_x[129] = c_Body_x[c_Size-1];
                        n_Body_y[129] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 130) begin
                        n_Body_x[130] = c_Body_x[129];
                        n_Body_y[130] = c_Body_y[129];
                    end else begin
                        n_Body_x[130] = c_Body_x[c_Size-1];
                        n_Body_y[130] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 131) begin
                        n_Body_x[131] = c_Body_x[130];
                        n_Body_y[131] = c_Body_y[130];
                    end else begin
                        n_Body_x[131] = c_Body_x[c_Size-1];
                        n_Body_y[131] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 132) begin
                        n_Body_x[132] = c_Body_x[131];
                        n_Body_y[132] = c_Body_y[131];
                    end else begin
                        n_Body_x[132] = c_Body_x[c_Size-1];
                        n_Body_y[132] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 133) begin
                        n_Body_x[133] = c_Body_x[132];
                        n_Body_y[133] = c_Body_y[132];
                    end else begin
                        n_Body_x[133] = c_Body_x[c_Size-1];
                        n_Body_y[133] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 134) begin
                        n_Body_x[134] = c_Body_x[133];
                        n_Body_y[134] = c_Body_y[133];
                    end else begin
                        n_Body_x[134] = c_Body_x[c_Size-1];
                        n_Body_y[134] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 135) begin
                        n_Body_x[135] = c_Body_x[134];
                        n_Body_y[135] = c_Body_y[134];
                    end else begin
                        n_Body_x[135] = c_Body_x[c_Size-1];
                        n_Body_y[135] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 136) begin
                        n_Body_x[136] = c_Body_x[135];
                        n_Body_y[136] = c_Body_y[135];
                    end else begin
                        n_Body_x[136] = c_Body_x[c_Size-1];
                        n_Body_y[136] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 137) begin
                        n_Body_x[137] = c_Body_x[136];
                        n_Body_y[137] = c_Body_y[136];
                    end else begin
                        n_Body_x[137] = c_Body_x[c_Size-1];
                        n_Body_y[137] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 138) begin
                        n_Body_x[138] = c_Body_x[137];
                        n_Body_y[138] = c_Body_y[137];
                    end else begin
                        n_Body_x[138] = c_Body_x[c_Size-1];
                        n_Body_y[138] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 139) begin
                        n_Body_x[139] = c_Body_x[138];
                        n_Body_y[139] = c_Body_y[138];
                    end else begin
                        n_Body_x[139] = c_Body_x[c_Size-1];
                        n_Body_y[139] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 140) begin
                        n_Body_x[140] = c_Body_x[139];
                        n_Body_y[140] = c_Body_y[139];
                    end else begin
                        n_Body_x[140] = c_Body_x[c_Size-1];
                        n_Body_y[140] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 141) begin
                        n_Body_x[141] = c_Body_x[140];
                        n_Body_y[141] = c_Body_y[140];
                    end else begin
                        n_Body_x[141] = c_Body_x[c_Size-1];
                        n_Body_y[141] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 142) begin
                        n_Body_x[142] = c_Body_x[141];
                        n_Body_y[142] = c_Body_y[141];
                    end else begin
                        n_Body_x[142] = c_Body_x[c_Size-1];
                        n_Body_y[142] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 143) begin
                        n_Body_x[143] = c_Body_x[142];
                        n_Body_y[143] = c_Body_y[142];
                    end else begin
                        n_Body_x[143] = c_Body_x[c_Size-1];
                        n_Body_y[143] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 144) begin
                        n_Body_x[144] = c_Body_x[143];
                        n_Body_y[144] = c_Body_y[143];
                    end else begin
                        n_Body_x[144] = c_Body_x[c_Size-1];
                        n_Body_y[144] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 145) begin
                        n_Body_x[145] = c_Body_x[144];
                        n_Body_y[145] = c_Body_y[144];
                    end else begin
                        n_Body_x[145] = c_Body_x[c_Size-1];
                        n_Body_y[145] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 146) begin
                        n_Body_x[146] = c_Body_x[145];
                        n_Body_y[146] = c_Body_y[145];
                    end else begin
                        n_Body_x[146] = c_Body_x[c_Size-1];
                        n_Body_y[146] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 147) begin
                        n_Body_x[147] = c_Body_x[146];
                        n_Body_y[147] = c_Body_y[146];
                    end else begin
                        n_Body_x[147] = c_Body_x[c_Size-1];
                        n_Body_y[147] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 148) begin
                        n_Body_x[148] = c_Body_x[147];
                        n_Body_y[148] = c_Body_y[147];
                    end else begin
                        n_Body_x[148] = c_Body_x[c_Size-1];
                        n_Body_y[148] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 149) begin
                        n_Body_x[149] = c_Body_x[148];
                        n_Body_y[149] = c_Body_y[148];
                    end else begin
                        n_Body_x[149] = c_Body_x[c_Size-1];
                        n_Body_y[149] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 150) begin
                        n_Body_x[150] = c_Body_x[149];
                        n_Body_y[150] = c_Body_y[149];
                    end else begin
                        n_Body_x[150] = c_Body_x[c_Size-1];
                        n_Body_y[150] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 151) begin
                        n_Body_x[151] = c_Body_x[150];
                        n_Body_y[151] = c_Body_y[150];
                    end else begin
                        n_Body_x[151] = c_Body_x[c_Size-1];
                        n_Body_y[151] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 152) begin
                        n_Body_x[152] = c_Body_x[151];
                        n_Body_y[152] = c_Body_y[151];
                    end else begin
                        n_Body_x[152] = c_Body_x[c_Size-1];
                        n_Body_y[152] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 153) begin
                        n_Body_x[153] = c_Body_x[152];
                        n_Body_y[153] = c_Body_y[152];
                    end else begin
                        n_Body_x[153] = c_Body_x[c_Size-1];
                        n_Body_y[153] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 154) begin
                        n_Body_x[154] = c_Body_x[153];
                        n_Body_y[154] = c_Body_y[153];
                    end else begin
                        n_Body_x[154] = c_Body_x[c_Size-1];
                        n_Body_y[154] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 155) begin
                        n_Body_x[155] = c_Body_x[154];
                        n_Body_y[155] = c_Body_y[154];
                    end else begin
                        n_Body_x[155] = c_Body_x[c_Size-1];
                        n_Body_y[155] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 156) begin
                        n_Body_x[156] = c_Body_x[155];
                        n_Body_y[156] = c_Body_y[155];
                    end else begin
                        n_Body_x[156] = c_Body_x[c_Size-1];
                        n_Body_y[156] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 157) begin
                        n_Body_x[157] = c_Body_x[156];
                        n_Body_y[157] = c_Body_y[156];
                    end else begin
                        n_Body_x[157] = c_Body_x[c_Size-1];
                        n_Body_y[157] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 158) begin
                        n_Body_x[158] = c_Body_x[157];
                        n_Body_y[158] = c_Body_y[157];
                    end else begin
                        n_Body_x[158] = c_Body_x[c_Size-1];
                        n_Body_y[158] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 159) begin
                        n_Body_x[159] = c_Body_x[158];
                        n_Body_y[159] = c_Body_y[158];
                    end else begin
                        n_Body_x[159] = c_Body_x[c_Size-1];
                        n_Body_y[159] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 160) begin
                        n_Body_x[160] = c_Body_x[159];
                        n_Body_y[160] = c_Body_y[159];
                    end else begin
                        n_Body_x[160] = c_Body_x[c_Size-1];
                        n_Body_y[160] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 161) begin
                        n_Body_x[161] = c_Body_x[160];
                        n_Body_y[161] = c_Body_y[160];
                    end else begin
                        n_Body_x[161] = c_Body_x[c_Size-1];
                        n_Body_y[161] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 162) begin
                        n_Body_x[162] = c_Body_x[161];
                        n_Body_y[162] = c_Body_y[161];
                    end else begin
                        n_Body_x[162] = c_Body_x[c_Size-1];
                        n_Body_y[162] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 163) begin
                        n_Body_x[163] = c_Body_x[162];
                        n_Body_y[163] = c_Body_y[162];
                    end else begin
                        n_Body_x[163] = c_Body_x[c_Size-1];
                        n_Body_y[163] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 164) begin
                        n_Body_x[164] = c_Body_x[163];
                        n_Body_y[164] = c_Body_y[163];
                    end else begin
                        n_Body_x[164] = c_Body_x[c_Size-1];
                        n_Body_y[164] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 165) begin
                        n_Body_x[165] = c_Body_x[164];
                        n_Body_y[165] = c_Body_y[164];
                    end else begin
                        n_Body_x[165] = c_Body_x[c_Size-1];
                        n_Body_y[165] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 166) begin
                        n_Body_x[166] = c_Body_x[165];
                        n_Body_y[166] = c_Body_y[165];
                    end else begin
                        n_Body_x[166] = c_Body_x[c_Size-1];
                        n_Body_y[166] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 167) begin
                        n_Body_x[167] = c_Body_x[166];
                        n_Body_y[167] = c_Body_y[166];
                    end else begin
                        n_Body_x[167] = c_Body_x[c_Size-1];
                        n_Body_y[167] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 168) begin
                        n_Body_x[168] = c_Body_x[167];
                        n_Body_y[168] = c_Body_y[167];
                    end else begin
                        n_Body_x[168] = c_Body_x[c_Size-1];
                        n_Body_y[168] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 169) begin
                        n_Body_x[169] = c_Body_x[168];
                        n_Body_y[169] = c_Body_y[168];
                    end else begin
                        n_Body_x[169] = c_Body_x[c_Size-1];
                        n_Body_y[169] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 170) begin
                        n_Body_x[170] = c_Body_x[169];
                        n_Body_y[170] = c_Body_y[169];
                    end else begin
                        n_Body_x[170] = c_Body_x[c_Size-1];
                        n_Body_y[170] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 171) begin
                        n_Body_x[171] = c_Body_x[170];
                        n_Body_y[171] = c_Body_y[170];
                    end else begin
                        n_Body_x[171] = c_Body_x[c_Size-1];
                        n_Body_y[171] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 172) begin
                        n_Body_x[172] = c_Body_x[171];
                        n_Body_y[172] = c_Body_y[171];
                    end else begin
                        n_Body_x[172] = c_Body_x[c_Size-1];
                        n_Body_y[172] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 173) begin
                        n_Body_x[173] = c_Body_x[172];
                        n_Body_y[173] = c_Body_y[172];
                    end else begin
                        n_Body_x[173] = c_Body_x[c_Size-1];
                        n_Body_y[173] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 174) begin
                        n_Body_x[174] = c_Body_x[173];
                        n_Body_y[174] = c_Body_y[173];
                    end else begin
                        n_Body_x[174] = c_Body_x[c_Size-1];
                        n_Body_y[174] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 175) begin
                        n_Body_x[175] = c_Body_x[174];
                        n_Body_y[175] = c_Body_y[174];
                    end else begin
                        n_Body_x[175] = c_Body_x[c_Size-1];
                        n_Body_y[175] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 176) begin
                        n_Body_x[176] = c_Body_x[175];
                        n_Body_y[176] = c_Body_y[175];
                    end else begin
                        n_Body_x[176] = c_Body_x[c_Size-1];
                        n_Body_y[176] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 177) begin
                        n_Body_x[177] = c_Body_x[176];
                        n_Body_y[177] = c_Body_y[176];
                    end else begin
                        n_Body_x[177] = c_Body_x[c_Size-1];
                        n_Body_y[177] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 178) begin
                        n_Body_x[178] = c_Body_x[177];
                        n_Body_y[178] = c_Body_y[177];
                    end else begin
                        n_Body_x[178] = c_Body_x[c_Size-1];
                        n_Body_y[178] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 179) begin
                        n_Body_x[179] = c_Body_x[178];
                        n_Body_y[179] = c_Body_y[178];
                    end else begin
                        n_Body_x[179] = c_Body_x[c_Size-1];
                        n_Body_y[179] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 180) begin
                        n_Body_x[180] = c_Body_x[179];
                        n_Body_y[180] = c_Body_y[179];
                    end else begin
                        n_Body_x[180] = c_Body_x[c_Size-1];
                        n_Body_y[180] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 181) begin
                        n_Body_x[181] = c_Body_x[180];
                        n_Body_y[181] = c_Body_y[180];
                    end else begin
                        n_Body_x[181] = c_Body_x[c_Size-1];
                        n_Body_y[181] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 182) begin
                        n_Body_x[182] = c_Body_x[181];
                        n_Body_y[182] = c_Body_y[181];
                    end else begin
                        n_Body_x[182] = c_Body_x[c_Size-1];
                        n_Body_y[182] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 183) begin
                        n_Body_x[183] = c_Body_x[182];
                        n_Body_y[183] = c_Body_y[182];
                    end else begin
                        n_Body_x[183] = c_Body_x[c_Size-1];
                        n_Body_y[183] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 184) begin
                        n_Body_x[184] = c_Body_x[183];
                        n_Body_y[184] = c_Body_y[183];
                    end else begin
                        n_Body_x[184] = c_Body_x[c_Size-1];
                        n_Body_y[184] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 185) begin
                        n_Body_x[185] = c_Body_x[184];
                        n_Body_y[185] = c_Body_y[184];
                    end else begin
                        n_Body_x[185] = c_Body_x[c_Size-1];
                        n_Body_y[185] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 186) begin
                        n_Body_x[186] = c_Body_x[185];
                        n_Body_y[186] = c_Body_y[185];
                    end else begin
                        n_Body_x[186] = c_Body_x[c_Size-1];
                        n_Body_y[186] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 187) begin
                        n_Body_x[187] = c_Body_x[186];
                        n_Body_y[187] = c_Body_y[186];
                    end else begin
                        n_Body_x[187] = c_Body_x[c_Size-1];
                        n_Body_y[187] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 188) begin
                        n_Body_x[188] = c_Body_x[187];
                        n_Body_y[188] = c_Body_y[187];
                    end else begin
                        n_Body_x[188] = c_Body_x[c_Size-1];
                        n_Body_y[188] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 189) begin
                        n_Body_x[189] = c_Body_x[188];
                        n_Body_y[189] = c_Body_y[188];
                    end else begin
                        n_Body_x[189] = c_Body_x[c_Size-1];
                        n_Body_y[189] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 190) begin
                        n_Body_x[190] = c_Body_x[189];
                        n_Body_y[190] = c_Body_y[189];
                    end else begin
                        n_Body_x[190] = c_Body_x[c_Size-1];
                        n_Body_y[190] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 191) begin
                        n_Body_x[191] = c_Body_x[190];
                        n_Body_y[191] = c_Body_y[190];
                    end else begin
                        n_Body_x[191] = c_Body_x[c_Size-1];
                        n_Body_y[191] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 192) begin
                        n_Body_x[192] = c_Body_x[191];
                        n_Body_y[192] = c_Body_y[191];
                    end else begin
                        n_Body_x[192] = c_Body_x[c_Size-1];
                        n_Body_y[192] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 193) begin
                        n_Body_x[193] = c_Body_x[192];
                        n_Body_y[193] = c_Body_y[192];
                    end else begin
                        n_Body_x[193] = c_Body_x[c_Size-1];
                        n_Body_y[193] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 194) begin
                        n_Body_x[194] = c_Body_x[193];
                        n_Body_y[194] = c_Body_y[193];
                    end else begin
                        n_Body_x[194] = c_Body_x[c_Size-1];
                        n_Body_y[194] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 195) begin
                        n_Body_x[195] = c_Body_x[194];
                        n_Body_y[195] = c_Body_y[194];
                    end else begin
                        n_Body_x[195] = c_Body_x[c_Size-1];
                        n_Body_y[195] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 196) begin
                        n_Body_x[196] = c_Body_x[195];
                        n_Body_y[196] = c_Body_y[195];
                    end else begin
                        n_Body_x[196] = c_Body_x[c_Size-1];
                        n_Body_y[196] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 197) begin
                        n_Body_x[197] = c_Body_x[196];
                        n_Body_y[197] = c_Body_y[196];
                    end else begin
                        n_Body_x[197] = c_Body_x[c_Size-1];
                        n_Body_y[197] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 198) begin
                        n_Body_x[198] = c_Body_x[197];
                        n_Body_y[198] = c_Body_y[197];
                    end else begin
                        n_Body_x[198] = c_Body_x[c_Size-1];
                        n_Body_y[198] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 199) begin
                        n_Body_x[199] = c_Body_x[198];
                        n_Body_y[199] = c_Body_y[198];
                    end else begin
                        n_Body_x[199] = c_Body_x[c_Size-1];
                        n_Body_y[199] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 200) begin
                        n_Body_x[200] = c_Body_x[199];
                        n_Body_y[200] = c_Body_y[199];
                    end else begin
                        n_Body_x[200] = c_Body_x[c_Size-1];
                        n_Body_y[200] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 201) begin
                        n_Body_x[201] = c_Body_x[200];
                        n_Body_y[201] = c_Body_y[200];
                    end else begin
                        n_Body_x[201] = c_Body_x[c_Size-1];
                        n_Body_y[201] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 202) begin
                        n_Body_x[202] = c_Body_x[201];
                        n_Body_y[202] = c_Body_y[201];
                    end else begin
                        n_Body_x[202] = c_Body_x[c_Size-1];
                        n_Body_y[202] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 203) begin
                        n_Body_x[203] = c_Body_x[202];
                        n_Body_y[203] = c_Body_y[202];
                    end else begin
                        n_Body_x[203] = c_Body_x[c_Size-1];
                        n_Body_y[203] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 204) begin
                        n_Body_x[204] = c_Body_x[203];
                        n_Body_y[204] = c_Body_y[203];
                    end else begin
                        n_Body_x[204] = c_Body_x[c_Size-1];
                        n_Body_y[204] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 205) begin
                        n_Body_x[205] = c_Body_x[204];
                        n_Body_y[205] = c_Body_y[204];
                    end else begin
                        n_Body_x[205] = c_Body_x[c_Size-1];
                        n_Body_y[205] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 206) begin
                        n_Body_x[206] = c_Body_x[205];
                        n_Body_y[206] = c_Body_y[205];
                    end else begin
                        n_Body_x[206] = c_Body_x[c_Size-1];
                        n_Body_y[206] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 207) begin
                        n_Body_x[207] = c_Body_x[206];
                        n_Body_y[207] = c_Body_y[206];
                    end else begin
                        n_Body_x[207] = c_Body_x[c_Size-1];
                        n_Body_y[207] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 208) begin
                        n_Body_x[208] = c_Body_x[207];
                        n_Body_y[208] = c_Body_y[207];
                    end else begin
                        n_Body_x[208] = c_Body_x[c_Size-1];
                        n_Body_y[208] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 209) begin
                        n_Body_x[209] = c_Body_x[208];
                        n_Body_y[209] = c_Body_y[208];
                    end else begin
                        n_Body_x[209] = c_Body_x[c_Size-1];
                        n_Body_y[209] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 210) begin
                        n_Body_x[210] = c_Body_x[209];
                        n_Body_y[210] = c_Body_y[209];
                    end else begin
                        n_Body_x[210] = c_Body_x[c_Size-1];
                        n_Body_y[210] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 211) begin
                        n_Body_x[211] = c_Body_x[210];
                        n_Body_y[211] = c_Body_y[210];
                    end else begin
                        n_Body_x[211] = c_Body_x[c_Size-1];
                        n_Body_y[211] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 212) begin
                        n_Body_x[212] = c_Body_x[211];
                        n_Body_y[212] = c_Body_y[211];
                    end else begin
                        n_Body_x[212] = c_Body_x[c_Size-1];
                        n_Body_y[212] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 213) begin
                        n_Body_x[213] = c_Body_x[212];
                        n_Body_y[213] = c_Body_y[212];
                    end else begin
                        n_Body_x[213] = c_Body_x[c_Size-1];
                        n_Body_y[213] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 214) begin
                        n_Body_x[214] = c_Body_x[213];
                        n_Body_y[214] = c_Body_y[213];
                    end else begin
                        n_Body_x[214] = c_Body_x[c_Size-1];
                        n_Body_y[214] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 215) begin
                        n_Body_x[215] = c_Body_x[214];
                        n_Body_y[215] = c_Body_y[214];
                    end else begin
                        n_Body_x[215] = c_Body_x[c_Size-1];
                        n_Body_y[215] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 216) begin
                        n_Body_x[216] = c_Body_x[215];
                        n_Body_y[216] = c_Body_y[215];
                    end else begin
                        n_Body_x[216] = c_Body_x[c_Size-1];
                        n_Body_y[216] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 217) begin
                        n_Body_x[217] = c_Body_x[216];
                        n_Body_y[217] = c_Body_y[216];
                    end else begin
                        n_Body_x[217] = c_Body_x[c_Size-1];
                        n_Body_y[217] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 218) begin
                        n_Body_x[218] = c_Body_x[217];
                        n_Body_y[218] = c_Body_y[217];
                    end else begin
                        n_Body_x[218] = c_Body_x[c_Size-1];
                        n_Body_y[218] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 219) begin
                        n_Body_x[219] = c_Body_x[218];
                        n_Body_y[219] = c_Body_y[218];
                    end else begin
                        n_Body_x[219] = c_Body_x[c_Size-1];
                        n_Body_y[219] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 220) begin
                        n_Body_x[220] = c_Body_x[219];
                        n_Body_y[220] = c_Body_y[219];
                    end else begin
                        n_Body_x[220] = c_Body_x[c_Size-1];
                        n_Body_y[220] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 221) begin
                        n_Body_x[221] = c_Body_x[220];
                        n_Body_y[221] = c_Body_y[220];
                    end else begin
                        n_Body_x[221] = c_Body_x[c_Size-1];
                        n_Body_y[221] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 222) begin
                        n_Body_x[222] = c_Body_x[221];
                        n_Body_y[222] = c_Body_y[221];
                    end else begin
                        n_Body_x[222] = c_Body_x[c_Size-1];
                        n_Body_y[222] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 223) begin
                        n_Body_x[223] = c_Body_x[222];
                        n_Body_y[223] = c_Body_y[222];
                    end else begin
                        n_Body_x[223] = c_Body_x[c_Size-1];
                        n_Body_y[223] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 224) begin
                        n_Body_x[224] = c_Body_x[223];
                        n_Body_y[224] = c_Body_y[223];
                    end else begin
                        n_Body_x[224] = c_Body_x[c_Size-1];
                        n_Body_y[224] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 225) begin
                        n_Body_x[225] = c_Body_x[224];
                        n_Body_y[225] = c_Body_y[224];
                    end else begin
                        n_Body_x[225] = c_Body_x[c_Size-1];
                        n_Body_y[225] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 226) begin
                        n_Body_x[226] = c_Body_x[225];
                        n_Body_y[226] = c_Body_y[225];
                    end else begin
                        n_Body_x[226] = c_Body_x[c_Size-1];
                        n_Body_y[226] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 227) begin
                        n_Body_x[227] = c_Body_x[226];
                        n_Body_y[227] = c_Body_y[226];
                    end else begin
                        n_Body_x[227] = c_Body_x[c_Size-1];
                        n_Body_y[227] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 228) begin
                        n_Body_x[228] = c_Body_x[227];
                        n_Body_y[228] = c_Body_y[227];
                    end else begin
                        n_Body_x[228] = c_Body_x[c_Size-1];
                        n_Body_y[228] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 229) begin
                        n_Body_x[229] = c_Body_x[228];
                        n_Body_y[229] = c_Body_y[228];
                    end else begin
                        n_Body_x[229] = c_Body_x[c_Size-1];
                        n_Body_y[229] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 230) begin
                        n_Body_x[230] = c_Body_x[229];
                        n_Body_y[230] = c_Body_y[229];
                    end else begin
                        n_Body_x[230] = c_Body_x[c_Size-1];
                        n_Body_y[230] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 231) begin
                        n_Body_x[231] = c_Body_x[230];
                        n_Body_y[231] = c_Body_y[230];
                    end else begin
                        n_Body_x[231] = c_Body_x[c_Size-1];
                        n_Body_y[231] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 232) begin
                        n_Body_x[232] = c_Body_x[231];
                        n_Body_y[232] = c_Body_y[231];
                    end else begin
                        n_Body_x[232] = c_Body_x[c_Size-1];
                        n_Body_y[232] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 233) begin
                        n_Body_x[233] = c_Body_x[232];
                        n_Body_y[233] = c_Body_y[232];
                    end else begin
                        n_Body_x[233] = c_Body_x[c_Size-1];
                        n_Body_y[233] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 234) begin
                        n_Body_x[234] = c_Body_x[233];
                        n_Body_y[234] = c_Body_y[233];
                    end else begin
                        n_Body_x[234] = c_Body_x[c_Size-1];
                        n_Body_y[234] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 235) begin
                        n_Body_x[235] = c_Body_x[234];
                        n_Body_y[235] = c_Body_y[234];
                    end else begin
                        n_Body_x[235] = c_Body_x[c_Size-1];
                        n_Body_y[235] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 236) begin
                        n_Body_x[236] = c_Body_x[235];
                        n_Body_y[236] = c_Body_y[235];
                    end else begin
                        n_Body_x[236] = c_Body_x[c_Size-1];
                        n_Body_y[236] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 237) begin
                        n_Body_x[237] = c_Body_x[236];
                        n_Body_y[237] = c_Body_y[236];
                    end else begin
                        n_Body_x[237] = c_Body_x[c_Size-1];
                        n_Body_y[237] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 238) begin
                        n_Body_x[238] = c_Body_x[237];
                        n_Body_y[238] = c_Body_y[237];
                    end else begin
                        n_Body_x[238] = c_Body_x[c_Size-1];
                        n_Body_y[238] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 239) begin
                        n_Body_x[239] = c_Body_x[238];
                        n_Body_y[239] = c_Body_y[238];
                    end else begin
                        n_Body_x[239] = c_Body_x[c_Size-1];
                        n_Body_y[239] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 240) begin
                        n_Body_x[240] = c_Body_x[239];
                        n_Body_y[240] = c_Body_y[239];
                    end else begin
                        n_Body_x[240] = c_Body_x[c_Size-1];
                        n_Body_y[240] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 241) begin
                        n_Body_x[241] = c_Body_x[240];
                        n_Body_y[241] = c_Body_y[240];
                    end else begin
                        n_Body_x[241] = c_Body_x[c_Size-1];
                        n_Body_y[241] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 242) begin
                        n_Body_x[242] = c_Body_x[241];
                        n_Body_y[242] = c_Body_y[241];
                    end else begin
                        n_Body_x[242] = c_Body_x[c_Size-1];
                        n_Body_y[242] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 243) begin
                        n_Body_x[243] = c_Body_x[242];
                        n_Body_y[243] = c_Body_y[242];
                    end else begin
                        n_Body_x[243] = c_Body_x[c_Size-1];
                        n_Body_y[243] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 244) begin
                        n_Body_x[244] = c_Body_x[243];
                        n_Body_y[244] = c_Body_y[243];
                    end else begin
                        n_Body_x[244] = c_Body_x[c_Size-1];
                        n_Body_y[244] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 245) begin
                        n_Body_x[245] = c_Body_x[244];
                        n_Body_y[245] = c_Body_y[244];
                    end else begin
                        n_Body_x[245] = c_Body_x[c_Size-1];
                        n_Body_y[245] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 246) begin
                        n_Body_x[246] = c_Body_x[245];
                        n_Body_y[246] = c_Body_y[245];
                    end else begin
                        n_Body_x[246] = c_Body_x[c_Size-1];
                        n_Body_y[246] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 247) begin
                        n_Body_x[247] = c_Body_x[246];
                        n_Body_y[247] = c_Body_y[246];
                    end else begin
                        n_Body_x[247] = c_Body_x[c_Size-1];
                        n_Body_y[247] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 248) begin
                        n_Body_x[248] = c_Body_x[247];
                        n_Body_y[248] = c_Body_y[247];
                    end else begin
                        n_Body_x[248] = c_Body_x[c_Size-1];
                        n_Body_y[248] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 249) begin
                        n_Body_x[249] = c_Body_x[248];
                        n_Body_y[249] = c_Body_y[248];
                    end else begin
                        n_Body_x[249] = c_Body_x[c_Size-1];
                        n_Body_y[249] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 250) begin
                        n_Body_x[250] = c_Body_x[249];
                        n_Body_y[250] = c_Body_y[249];
                    end else begin
                        n_Body_x[250] = c_Body_x[c_Size-1];
                        n_Body_y[250] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 251) begin
                        n_Body_x[251] = c_Body_x[250];
                        n_Body_y[251] = c_Body_y[250];
                    end else begin
                        n_Body_x[251] = c_Body_x[c_Size-1];
                        n_Body_y[251] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 252) begin
                        n_Body_x[252] = c_Body_x[251];
                        n_Body_y[252] = c_Body_y[251];
                    end else begin
                        n_Body_x[252] = c_Body_x[c_Size-1];
                        n_Body_y[252] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 253) begin
                        n_Body_x[253] = c_Body_x[252];
                        n_Body_y[253] = c_Body_y[252];
                    end else begin
                        n_Body_x[253] = c_Body_x[c_Size-1];
                        n_Body_y[253] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 254) begin
                        n_Body_x[254] = c_Body_x[253];
                        n_Body_y[254] = c_Body_y[253];
                    end else begin
                        n_Body_x[254] = c_Body_x[c_Size-1];
                        n_Body_y[254] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 255) begin
                        n_Body_x[255] = c_Body_x[254];
                        n_Body_y[255] = c_Body_y[254];
                    end else begin
                        n_Body_x[255] = c_Body_x[c_Size-1];
                        n_Body_y[255] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 256) begin
                        n_Body_x[256] = c_Body_x[255];
                        n_Body_y[256] = c_Body_y[255];
                    end else begin
                        n_Body_x[256] = c_Body_x[c_Size-1];
                        n_Body_y[256] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 257) begin
                        n_Body_x[257] = c_Body_x[256];
                        n_Body_y[257] = c_Body_y[256];
                    end else begin
                        n_Body_x[257] = c_Body_x[c_Size-1];
                        n_Body_y[257] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 258) begin
                        n_Body_x[258] = c_Body_x[257];
                        n_Body_y[258] = c_Body_y[257];
                    end else begin
                        n_Body_x[258] = c_Body_x[c_Size-1];
                        n_Body_y[258] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 259) begin
                        n_Body_x[259] = c_Body_x[258];
                        n_Body_y[259] = c_Body_y[258];
                    end else begin
                        n_Body_x[259] = c_Body_x[c_Size-1];
                        n_Body_y[259] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 260) begin
                        n_Body_x[260] = c_Body_x[259];
                        n_Body_y[260] = c_Body_y[259];
                    end else begin
                        n_Body_x[260] = c_Body_x[c_Size-1];
                        n_Body_y[260] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 261) begin
                        n_Body_x[261] = c_Body_x[260];
                        n_Body_y[261] = c_Body_y[260];
                    end else begin
                        n_Body_x[261] = c_Body_x[c_Size-1];
                        n_Body_y[261] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 262) begin
                        n_Body_x[262] = c_Body_x[261];
                        n_Body_y[262] = c_Body_y[261];
                    end else begin
                        n_Body_x[262] = c_Body_x[c_Size-1];
                        n_Body_y[262] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 263) begin
                        n_Body_x[263] = c_Body_x[262];
                        n_Body_y[263] = c_Body_y[262];
                    end else begin
                        n_Body_x[263] = c_Body_x[c_Size-1];
                        n_Body_y[263] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 264) begin
                        n_Body_x[264] = c_Body_x[263];
                        n_Body_y[264] = c_Body_y[263];
                    end else begin
                        n_Body_x[264] = c_Body_x[c_Size-1];
                        n_Body_y[264] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 265) begin
                        n_Body_x[265] = c_Body_x[264];
                        n_Body_y[265] = c_Body_y[264];
                    end else begin
                        n_Body_x[265] = c_Body_x[c_Size-1];
                        n_Body_y[265] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 266) begin
                        n_Body_x[266] = c_Body_x[265];
                        n_Body_y[266] = c_Body_y[265];
                    end else begin
                        n_Body_x[266] = c_Body_x[c_Size-1];
                        n_Body_y[266] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 267) begin
                        n_Body_x[267] = c_Body_x[266];
                        n_Body_y[267] = c_Body_y[266];
                    end else begin
                        n_Body_x[267] = c_Body_x[c_Size-1];
                        n_Body_y[267] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 268) begin
                        n_Body_x[268] = c_Body_x[267];
                        n_Body_y[268] = c_Body_y[267];
                    end else begin
                        n_Body_x[268] = c_Body_x[c_Size-1];
                        n_Body_y[268] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 269) begin
                        n_Body_x[269] = c_Body_x[268];
                        n_Body_y[269] = c_Body_y[268];
                    end else begin
                        n_Body_x[269] = c_Body_x[c_Size-1];
                        n_Body_y[269] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 270) begin
                        n_Body_x[270] = c_Body_x[269];
                        n_Body_y[270] = c_Body_y[269];
                    end else begin
                        n_Body_x[270] = c_Body_x[c_Size-1];
                        n_Body_y[270] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 271) begin
                        n_Body_x[271] = c_Body_x[270];
                        n_Body_y[271] = c_Body_y[270];
                    end else begin
                        n_Body_x[271] = c_Body_x[c_Size-1];
                        n_Body_y[271] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 272) begin
                        n_Body_x[272] = c_Body_x[271];
                        n_Body_y[272] = c_Body_y[271];
                    end else begin
                        n_Body_x[272] = c_Body_x[c_Size-1];
                        n_Body_y[272] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 273) begin
                        n_Body_x[273] = c_Body_x[272];
                        n_Body_y[273] = c_Body_y[272];
                    end else begin
                        n_Body_x[273] = c_Body_x[c_Size-1];
                        n_Body_y[273] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 274) begin
                        n_Body_x[274] = c_Body_x[273];
                        n_Body_y[274] = c_Body_y[273];
                    end else begin
                        n_Body_x[274] = c_Body_x[c_Size-1];
                        n_Body_y[274] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 275) begin
                        n_Body_x[275] = c_Body_x[274];
                        n_Body_y[275] = c_Body_y[274];
                    end else begin
                        n_Body_x[275] = c_Body_x[c_Size-1];
                        n_Body_y[275] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 276) begin
                        n_Body_x[276] = c_Body_x[275];
                        n_Body_y[276] = c_Body_y[275];
                    end else begin
                        n_Body_x[276] = c_Body_x[c_Size-1];
                        n_Body_y[276] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 277) begin
                        n_Body_x[277] = c_Body_x[276];
                        n_Body_y[277] = c_Body_y[276];
                    end else begin
                        n_Body_x[277] = c_Body_x[c_Size-1];
                        n_Body_y[277] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 278) begin
                        n_Body_x[278] = c_Body_x[277];
                        n_Body_y[278] = c_Body_y[277];
                    end else begin
                        n_Body_x[278] = c_Body_x[c_Size-1];
                        n_Body_y[278] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 279) begin
                        n_Body_x[279] = c_Body_x[278];
                        n_Body_y[279] = c_Body_y[278];
                    end else begin
                        n_Body_x[279] = c_Body_x[c_Size-1];
                        n_Body_y[279] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 280) begin
                        n_Body_x[280] = c_Body_x[279];
                        n_Body_y[280] = c_Body_y[279];
                    end else begin
                        n_Body_x[280] = c_Body_x[c_Size-1];
                        n_Body_y[280] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 281) begin
                        n_Body_x[281] = c_Body_x[280];
                        n_Body_y[281] = c_Body_y[280];
                    end else begin
                        n_Body_x[281] = c_Body_x[c_Size-1];
                        n_Body_y[281] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 282) begin
                        n_Body_x[282] = c_Body_x[281];
                        n_Body_y[282] = c_Body_y[281];
                    end else begin
                        n_Body_x[282] = c_Body_x[c_Size-1];
                        n_Body_y[282] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 283) begin
                        n_Body_x[283] = c_Body_x[282];
                        n_Body_y[283] = c_Body_y[282];
                    end else begin
                        n_Body_x[283] = c_Body_x[c_Size-1];
                        n_Body_y[283] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 284) begin
                        n_Body_x[284] = c_Body_x[283];
                        n_Body_y[284] = c_Body_y[283];
                    end else begin
                        n_Body_x[284] = c_Body_x[c_Size-1];
                        n_Body_y[284] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 285) begin
                        n_Body_x[285] = c_Body_x[284];
                        n_Body_y[285] = c_Body_y[284];
                    end else begin
                        n_Body_x[285] = c_Body_x[c_Size-1];
                        n_Body_y[285] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 286) begin
                        n_Body_x[286] = c_Body_x[285];
                        n_Body_y[286] = c_Body_y[285];
                    end else begin
                        n_Body_x[286] = c_Body_x[c_Size-1];
                        n_Body_y[286] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 287) begin
                        n_Body_x[287] = c_Body_x[286];
                        n_Body_y[287] = c_Body_y[286];
                    end else begin
                        n_Body_x[287] = c_Body_x[c_Size-1];
                        n_Body_y[287] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 288) begin
                        n_Body_x[288] = c_Body_x[287];
                        n_Body_y[288] = c_Body_y[287];
                    end else begin
                        n_Body_x[288] = c_Body_x[c_Size-1];
                        n_Body_y[288] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 289) begin
                        n_Body_x[289] = c_Body_x[288];
                        n_Body_y[289] = c_Body_y[288];
                    end else begin
                        n_Body_x[289] = c_Body_x[c_Size-1];
                        n_Body_y[289] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 290) begin
                        n_Body_x[290] = c_Body_x[289];
                        n_Body_y[290] = c_Body_y[289];
                    end else begin
                        n_Body_x[290] = c_Body_x[c_Size-1];
                        n_Body_y[290] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 291) begin
                        n_Body_x[291] = c_Body_x[290];
                        n_Body_y[291] = c_Body_y[290];
                    end else begin
                        n_Body_x[291] = c_Body_x[c_Size-1];
                        n_Body_y[291] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 292) begin
                        n_Body_x[292] = c_Body_x[291];
                        n_Body_y[292] = c_Body_y[291];
                    end else begin
                        n_Body_x[292] = c_Body_x[c_Size-1];
                        n_Body_y[292] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 293) begin
                        n_Body_x[293] = c_Body_x[292];
                        n_Body_y[293] = c_Body_y[292];
                    end else begin
                        n_Body_x[293] = c_Body_x[c_Size-1];
                        n_Body_y[293] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 294) begin
                        n_Body_x[294] = c_Body_x[293];
                        n_Body_y[294] = c_Body_y[293];
                    end else begin
                        n_Body_x[294] = c_Body_x[c_Size-1];
                        n_Body_y[294] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 295) begin
                        n_Body_x[295] = c_Body_x[294];
                        n_Body_y[295] = c_Body_y[294];
                    end else begin
                        n_Body_x[295] = c_Body_x[c_Size-1];
                        n_Body_y[295] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 296) begin
                        n_Body_x[296] = c_Body_x[295];
                        n_Body_y[296] = c_Body_y[295];
                    end else begin
                        n_Body_x[296] = c_Body_x[c_Size-1];
                        n_Body_y[296] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 297) begin
                        n_Body_x[297] = c_Body_x[296];
                        n_Body_y[297] = c_Body_y[296];
                    end else begin
                        n_Body_x[297] = c_Body_x[c_Size-1];
                        n_Body_y[297] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 298) begin
                        n_Body_x[298] = c_Body_x[297];
                        n_Body_y[298] = c_Body_y[297];
                    end else begin
                        n_Body_x[298] = c_Body_x[c_Size-1];
                        n_Body_y[298] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 299) begin
                        n_Body_x[299] = c_Body_x[298];
                        n_Body_y[299] = c_Body_y[298];
                    end else begin
                        n_Body_x[299] = c_Body_x[c_Size-1];
                        n_Body_y[299] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 300) begin
                        n_Body_x[300] = c_Body_x[299];
                        n_Body_y[300] = c_Body_y[299];
                    end else begin
                        n_Body_x[300] = c_Body_x[c_Size-1];
                        n_Body_y[300] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 301) begin
                        n_Body_x[301] = c_Body_x[300];
                        n_Body_y[301] = c_Body_y[300];
                    end else begin
                        n_Body_x[301] = c_Body_x[c_Size-1];
                        n_Body_y[301] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 302) begin
                        n_Body_x[302] = c_Body_x[301];
                        n_Body_y[302] = c_Body_y[301];
                    end else begin
                        n_Body_x[302] = c_Body_x[c_Size-1];
                        n_Body_y[302] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 303) begin
                        n_Body_x[303] = c_Body_x[302];
                        n_Body_y[303] = c_Body_y[302];
                    end else begin
                        n_Body_x[303] = c_Body_x[c_Size-1];
                        n_Body_y[303] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 304) begin
                        n_Body_x[304] = c_Body_x[303];
                        n_Body_y[304] = c_Body_y[303];
                    end else begin
                        n_Body_x[304] = c_Body_x[c_Size-1];
                        n_Body_y[304] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 305) begin
                        n_Body_x[305] = c_Body_x[304];
                        n_Body_y[305] = c_Body_y[304];
                    end else begin
                        n_Body_x[305] = c_Body_x[c_Size-1];
                        n_Body_y[305] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 306) begin
                        n_Body_x[306] = c_Body_x[305];
                        n_Body_y[306] = c_Body_y[305];
                    end else begin
                        n_Body_x[306] = c_Body_x[c_Size-1];
                        n_Body_y[306] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 307) begin
                        n_Body_x[307] = c_Body_x[306];
                        n_Body_y[307] = c_Body_y[306];
                    end else begin
                        n_Body_x[307] = c_Body_x[c_Size-1];
                        n_Body_y[307] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 308) begin
                        n_Body_x[308] = c_Body_x[307];
                        n_Body_y[308] = c_Body_y[307];
                    end else begin
                        n_Body_x[308] = c_Body_x[c_Size-1];
                        n_Body_y[308] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 309) begin
                        n_Body_x[309] = c_Body_x[308];
                        n_Body_y[309] = c_Body_y[308];
                    end else begin
                        n_Body_x[309] = c_Body_x[c_Size-1];
                        n_Body_y[309] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 310) begin
                        n_Body_x[310] = c_Body_x[309];
                        n_Body_y[310] = c_Body_y[309];
                    end else begin
                        n_Body_x[310] = c_Body_x[c_Size-1];
                        n_Body_y[310] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 311) begin
                        n_Body_x[311] = c_Body_x[310];
                        n_Body_y[311] = c_Body_y[310];
                    end else begin
                        n_Body_x[311] = c_Body_x[c_Size-1];
                        n_Body_y[311] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 312) begin
                        n_Body_x[312] = c_Body_x[311];
                        n_Body_y[312] = c_Body_y[311];
                    end else begin
                        n_Body_x[312] = c_Body_x[c_Size-1];
                        n_Body_y[312] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 313) begin
                        n_Body_x[313] = c_Body_x[312];
                        n_Body_y[313] = c_Body_y[312];
                    end else begin
                        n_Body_x[313] = c_Body_x[c_Size-1];
                        n_Body_y[313] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 314) begin
                        n_Body_x[314] = c_Body_x[313];
                        n_Body_y[314] = c_Body_y[313];
                    end else begin
                        n_Body_x[314] = c_Body_x[c_Size-1];
                        n_Body_y[314] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 315) begin
                        n_Body_x[315] = c_Body_x[314];
                        n_Body_y[315] = c_Body_y[314];
                    end else begin
                        n_Body_x[315] = c_Body_x[c_Size-1];
                        n_Body_y[315] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 316) begin
                        n_Body_x[316] = c_Body_x[315];
                        n_Body_y[316] = c_Body_y[315];
                    end else begin
                        n_Body_x[316] = c_Body_x[c_Size-1];
                        n_Body_y[316] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 317) begin
                        n_Body_x[317] = c_Body_x[316];
                        n_Body_y[317] = c_Body_y[316];
                    end else begin
                        n_Body_x[317] = c_Body_x[c_Size-1];
                        n_Body_y[317] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 318) begin
                        n_Body_x[318] = c_Body_x[317];
                        n_Body_y[318] = c_Body_y[317];
                    end else begin
                        n_Body_x[318] = c_Body_x[c_Size-1];
                        n_Body_y[318] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 319) begin
                        n_Body_x[319] = c_Body_x[318];
                        n_Body_y[319] = c_Body_y[318];
                    end else begin
                        n_Body_x[319] = c_Body_x[c_Size-1];
                        n_Body_y[319] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 320) begin
                        n_Body_x[320] = c_Body_x[319];
                        n_Body_y[320] = c_Body_y[319];
                    end else begin
                        n_Body_x[320] = c_Body_x[c_Size-1];
                        n_Body_y[320] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 321) begin
                        n_Body_x[321] = c_Body_x[320];
                        n_Body_y[321] = c_Body_y[320];
                    end else begin
                        n_Body_x[321] = c_Body_x[c_Size-1];
                        n_Body_y[321] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 322) begin
                        n_Body_x[322] = c_Body_x[321];
                        n_Body_y[322] = c_Body_y[321];
                    end else begin
                        n_Body_x[322] = c_Body_x[c_Size-1];
                        n_Body_y[322] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 323) begin
                        n_Body_x[323] = c_Body_x[322];
                        n_Body_y[323] = c_Body_y[322];
                    end else begin
                        n_Body_x[323] = c_Body_x[c_Size-1];
                        n_Body_y[323] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 324) begin
                        n_Body_x[324] = c_Body_x[323];
                        n_Body_y[324] = c_Body_y[323];
                    end else begin
                        n_Body_x[324] = c_Body_x[c_Size-1];
                        n_Body_y[324] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 325) begin
                        n_Body_x[325] = c_Body_x[324];
                        n_Body_y[325] = c_Body_y[324];
                    end else begin
                        n_Body_x[325] = c_Body_x[c_Size-1];
                        n_Body_y[325] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 326) begin
                        n_Body_x[326] = c_Body_x[325];
                        n_Body_y[326] = c_Body_y[325];
                    end else begin
                        n_Body_x[326] = c_Body_x[c_Size-1];
                        n_Body_y[326] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 327) begin
                        n_Body_x[327] = c_Body_x[326];
                        n_Body_y[327] = c_Body_y[326];
                    end else begin
                        n_Body_x[327] = c_Body_x[c_Size-1];
                        n_Body_y[327] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 328) begin
                        n_Body_x[328] = c_Body_x[327];
                        n_Body_y[328] = c_Body_y[327];
                    end else begin
                        n_Body_x[328] = c_Body_x[c_Size-1];
                        n_Body_y[328] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 329) begin
                        n_Body_x[329] = c_Body_x[328];
                        n_Body_y[329] = c_Body_y[328];
                    end else begin
                        n_Body_x[329] = c_Body_x[c_Size-1];
                        n_Body_y[329] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 330) begin
                        n_Body_x[330] = c_Body_x[329];
                        n_Body_y[330] = c_Body_y[329];
                    end else begin
                        n_Body_x[330] = c_Body_x[c_Size-1];
                        n_Body_y[330] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 331) begin
                        n_Body_x[331] = c_Body_x[330];
                        n_Body_y[331] = c_Body_y[330];
                    end else begin
                        n_Body_x[331] = c_Body_x[c_Size-1];
                        n_Body_y[331] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 332) begin
                        n_Body_x[332] = c_Body_x[331];
                        n_Body_y[332] = c_Body_y[331];
                    end else begin
                        n_Body_x[332] = c_Body_x[c_Size-1];
                        n_Body_y[332] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 333) begin
                        n_Body_x[333] = c_Body_x[332];
                        n_Body_y[333] = c_Body_y[332];
                    end else begin
                        n_Body_x[333] = c_Body_x[c_Size-1];
                        n_Body_y[333] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 334) begin
                        n_Body_x[334] = c_Body_x[333];
                        n_Body_y[334] = c_Body_y[333];
                    end else begin
                        n_Body_x[334] = c_Body_x[c_Size-1];
                        n_Body_y[334] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 335) begin
                        n_Body_x[335] = c_Body_x[334];
                        n_Body_y[335] = c_Body_y[334];
                    end else begin
                        n_Body_x[335] = c_Body_x[c_Size-1];
                        n_Body_y[335] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 336) begin
                        n_Body_x[336] = c_Body_x[335];
                        n_Body_y[336] = c_Body_y[335];
                    end else begin
                        n_Body_x[336] = c_Body_x[c_Size-1];
                        n_Body_y[336] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 337) begin
                        n_Body_x[337] = c_Body_x[336];
                        n_Body_y[337] = c_Body_y[336];
                    end else begin
                        n_Body_x[337] = c_Body_x[c_Size-1];
                        n_Body_y[337] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 338) begin
                        n_Body_x[338] = c_Body_x[337];
                        n_Body_y[338] = c_Body_y[337];
                    end else begin
                        n_Body_x[338] = c_Body_x[c_Size-1];
                        n_Body_y[338] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 339) begin
                        n_Body_x[339] = c_Body_x[338];
                        n_Body_y[339] = c_Body_y[338];
                    end else begin
                        n_Body_x[339] = c_Body_x[c_Size-1];
                        n_Body_y[339] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 340) begin
                        n_Body_x[340] = c_Body_x[339];
                        n_Body_y[340] = c_Body_y[339];
                    end else begin
                        n_Body_x[340] = c_Body_x[c_Size-1];
                        n_Body_y[340] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 341) begin
                        n_Body_x[341] = c_Body_x[340];
                        n_Body_y[341] = c_Body_y[340];
                    end else begin
                        n_Body_x[341] = c_Body_x[c_Size-1];
                        n_Body_y[341] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 342) begin
                        n_Body_x[342] = c_Body_x[341];
                        n_Body_y[342] = c_Body_y[341];
                    end else begin
                        n_Body_x[342] = c_Body_x[c_Size-1];
                        n_Body_y[342] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 343) begin
                        n_Body_x[343] = c_Body_x[342];
                        n_Body_y[343] = c_Body_y[342];
                    end else begin
                        n_Body_x[343] = c_Body_x[c_Size-1];
                        n_Body_y[343] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 344) begin
                        n_Body_x[344] = c_Body_x[343];
                        n_Body_y[344] = c_Body_y[343];
                    end else begin
                        n_Body_x[344] = c_Body_x[c_Size-1];
                        n_Body_y[344] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 345) begin
                        n_Body_x[345] = c_Body_x[344];
                        n_Body_y[345] = c_Body_y[344];
                    end else begin
                        n_Body_x[345] = c_Body_x[c_Size-1];
                        n_Body_y[345] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 346) begin
                        n_Body_x[346] = c_Body_x[345];
                        n_Body_y[346] = c_Body_y[345];
                    end else begin
                        n_Body_x[346] = c_Body_x[c_Size-1];
                        n_Body_y[346] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 347) begin
                        n_Body_x[347] = c_Body_x[346];
                        n_Body_y[347] = c_Body_y[346];
                    end else begin
                        n_Body_x[347] = c_Body_x[c_Size-1];
                        n_Body_y[347] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 348) begin
                        n_Body_x[348] = c_Body_x[347];
                        n_Body_y[348] = c_Body_y[347];
                    end else begin
                        n_Body_x[348] = c_Body_x[c_Size-1];
                        n_Body_y[348] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 349) begin
                        n_Body_x[349] = c_Body_x[348];
                        n_Body_y[349] = c_Body_y[348];
                    end else begin
                        n_Body_x[349] = c_Body_x[c_Size-1];
                        n_Body_y[349] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 350) begin
                        n_Body_x[350] = c_Body_x[349];
                        n_Body_y[350] = c_Body_y[349];
                    end else begin
                        n_Body_x[350] = c_Body_x[c_Size-1];
                        n_Body_y[350] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 351) begin
                        n_Body_x[351] = c_Body_x[350];
                        n_Body_y[351] = c_Body_y[350];
                    end else begin
                        n_Body_x[351] = c_Body_x[c_Size-1];
                        n_Body_y[351] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 352) begin
                        n_Body_x[352] = c_Body_x[351];
                        n_Body_y[352] = c_Body_y[351];
                    end else begin
                        n_Body_x[352] = c_Body_x[c_Size-1];
                        n_Body_y[352] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 353) begin
                        n_Body_x[353] = c_Body_x[352];
                        n_Body_y[353] = c_Body_y[352];
                    end else begin
                        n_Body_x[353] = c_Body_x[c_Size-1];
                        n_Body_y[353] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 354) begin
                        n_Body_x[354] = c_Body_x[353];
                        n_Body_y[354] = c_Body_y[353];
                    end else begin
                        n_Body_x[354] = c_Body_x[c_Size-1];
                        n_Body_y[354] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 355) begin
                        n_Body_x[355] = c_Body_x[354];
                        n_Body_y[355] = c_Body_y[354];
                    end else begin
                        n_Body_x[355] = c_Body_x[c_Size-1];
                        n_Body_y[355] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 356) begin
                        n_Body_x[356] = c_Body_x[355];
                        n_Body_y[356] = c_Body_y[355];
                    end else begin
                        n_Body_x[356] = c_Body_x[c_Size-1];
                        n_Body_y[356] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 357) begin
                        n_Body_x[357] = c_Body_x[356];
                        n_Body_y[357] = c_Body_y[356];
                    end else begin
                        n_Body_x[357] = c_Body_x[c_Size-1];
                        n_Body_y[357] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 358) begin
                        n_Body_x[358] = c_Body_x[357];
                        n_Body_y[358] = c_Body_y[357];
                    end else begin
                        n_Body_x[358] = c_Body_x[c_Size-1];
                        n_Body_y[358] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 359) begin
                        n_Body_x[359] = c_Body_x[358];
                        n_Body_y[359] = c_Body_y[358];
                    end else begin
                        n_Body_x[359] = c_Body_x[c_Size-1];
                        n_Body_y[359] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 360) begin
                        n_Body_x[360] = c_Body_x[359];
                        n_Body_y[360] = c_Body_y[359];
                    end else begin
                        n_Body_x[360] = c_Body_x[c_Size-1];
                        n_Body_y[360] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 361) begin
                        n_Body_x[361] = c_Body_x[360];
                        n_Body_y[361] = c_Body_y[360];
                    end else begin
                        n_Body_x[361] = c_Body_x[c_Size-1];
                        n_Body_y[361] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 362) begin
                        n_Body_x[362] = c_Body_x[361];
                        n_Body_y[362] = c_Body_y[361];
                    end else begin
                        n_Body_x[362] = c_Body_x[c_Size-1];
                        n_Body_y[362] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 363) begin
                        n_Body_x[363] = c_Body_x[362];
                        n_Body_y[363] = c_Body_y[362];
                    end else begin
                        n_Body_x[363] = c_Body_x[c_Size-1];
                        n_Body_y[363] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 364) begin
                        n_Body_x[364] = c_Body_x[363];
                        n_Body_y[364] = c_Body_y[363];
                    end else begin
                        n_Body_x[364] = c_Body_x[c_Size-1];
                        n_Body_y[364] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 365) begin
                        n_Body_x[365] = c_Body_x[364];
                        n_Body_y[365] = c_Body_y[364];
                    end else begin
                        n_Body_x[365] = c_Body_x[c_Size-1];
                        n_Body_y[365] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 366) begin
                        n_Body_x[366] = c_Body_x[365];
                        n_Body_y[366] = c_Body_y[365];
                    end else begin
                        n_Body_x[366] = c_Body_x[c_Size-1];
                        n_Body_y[366] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 367) begin
                        n_Body_x[367] = c_Body_x[366];
                        n_Body_y[367] = c_Body_y[366];
                    end else begin
                        n_Body_x[367] = c_Body_x[c_Size-1];
                        n_Body_y[367] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 368) begin
                        n_Body_x[368] = c_Body_x[367];
                        n_Body_y[368] = c_Body_y[367];
                    end else begin
                        n_Body_x[368] = c_Body_x[c_Size-1];
                        n_Body_y[368] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 369) begin
                        n_Body_x[369] = c_Body_x[368];
                        n_Body_y[369] = c_Body_y[368];
                    end else begin
                        n_Body_x[369] = c_Body_x[c_Size-1];
                        n_Body_y[369] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 370) begin
                        n_Body_x[370] = c_Body_x[369];
                        n_Body_y[370] = c_Body_y[369];
                    end else begin
                        n_Body_x[370] = c_Body_x[c_Size-1];
                        n_Body_y[370] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 371) begin
                        n_Body_x[371] = c_Body_x[370];
                        n_Body_y[371] = c_Body_y[370];
                    end else begin
                        n_Body_x[371] = c_Body_x[c_Size-1];
                        n_Body_y[371] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 372) begin
                        n_Body_x[372] = c_Body_x[371];
                        n_Body_y[372] = c_Body_y[371];
                    end else begin
                        n_Body_x[372] = c_Body_x[c_Size-1];
                        n_Body_y[372] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 373) begin
                        n_Body_x[373] = c_Body_x[372];
                        n_Body_y[373] = c_Body_y[372];
                    end else begin
                        n_Body_x[373] = c_Body_x[c_Size-1];
                        n_Body_y[373] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 374) begin
                        n_Body_x[374] = c_Body_x[373];
                        n_Body_y[374] = c_Body_y[373];
                    end else begin
                        n_Body_x[374] = c_Body_x[c_Size-1];
                        n_Body_y[374] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 375) begin
                        n_Body_x[375] = c_Body_x[374];
                        n_Body_y[375] = c_Body_y[374];
                    end else begin
                        n_Body_x[375] = c_Body_x[c_Size-1];
                        n_Body_y[375] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 376) begin
                        n_Body_x[376] = c_Body_x[375];
                        n_Body_y[376] = c_Body_y[375];
                    end else begin
                        n_Body_x[376] = c_Body_x[c_Size-1];
                        n_Body_y[376] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 377) begin
                        n_Body_x[377] = c_Body_x[376];
                        n_Body_y[377] = c_Body_y[376];
                    end else begin
                        n_Body_x[377] = c_Body_x[c_Size-1];
                        n_Body_y[377] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 378) begin
                        n_Body_x[378] = c_Body_x[377];
                        n_Body_y[378] = c_Body_y[377];
                    end else begin
                        n_Body_x[378] = c_Body_x[c_Size-1];
                        n_Body_y[378] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 379) begin
                        n_Body_x[379] = c_Body_x[378];
                        n_Body_y[379] = c_Body_y[378];
                    end else begin
                        n_Body_x[379] = c_Body_x[c_Size-1];
                        n_Body_y[379] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 380) begin
                        n_Body_x[380] = c_Body_x[379];
                        n_Body_y[380] = c_Body_y[379];
                    end else begin
                        n_Body_x[380] = c_Body_x[c_Size-1];
                        n_Body_y[380] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 381) begin
                        n_Body_x[381] = c_Body_x[380];
                        n_Body_y[381] = c_Body_y[380];
                    end else begin
                        n_Body_x[381] = c_Body_x[c_Size-1];
                        n_Body_y[381] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 382) begin
                        n_Body_x[382] = c_Body_x[381];
                        n_Body_y[382] = c_Body_y[381];
                    end else begin
                        n_Body_x[382] = c_Body_x[c_Size-1];
                        n_Body_y[382] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 383) begin
                        n_Body_x[383] = c_Body_x[382];
                        n_Body_y[383] = c_Body_y[382];
                    end else begin
                        n_Body_x[383] = c_Body_x[c_Size-1];
                        n_Body_y[383] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 384) begin
                        n_Body_x[384] = c_Body_x[383];
                        n_Body_y[384] = c_Body_y[383];
                    end else begin
                        n_Body_x[384] = c_Body_x[c_Size-1];
                        n_Body_y[384] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 385) begin
                        n_Body_x[385] = c_Body_x[384];
                        n_Body_y[385] = c_Body_y[384];
                    end else begin
                        n_Body_x[385] = c_Body_x[c_Size-1];
                        n_Body_y[385] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 386) begin
                        n_Body_x[386] = c_Body_x[385];
                        n_Body_y[386] = c_Body_y[385];
                    end else begin
                        n_Body_x[386] = c_Body_x[c_Size-1];
                        n_Body_y[386] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 387) begin
                        n_Body_x[387] = c_Body_x[386];
                        n_Body_y[387] = c_Body_y[386];
                    end else begin
                        n_Body_x[387] = c_Body_x[c_Size-1];
                        n_Body_y[387] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 388) begin
                        n_Body_x[388] = c_Body_x[387];
                        n_Body_y[388] = c_Body_y[387];
                    end else begin
                        n_Body_x[388] = c_Body_x[c_Size-1];
                        n_Body_y[388] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 389) begin
                        n_Body_x[389] = c_Body_x[388];
                        n_Body_y[389] = c_Body_y[388];
                    end else begin
                        n_Body_x[389] = c_Body_x[c_Size-1];
                        n_Body_y[389] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 390) begin
                        n_Body_x[390] = c_Body_x[389];
                        n_Body_y[390] = c_Body_y[389];
                    end else begin
                        n_Body_x[390] = c_Body_x[c_Size-1];
                        n_Body_y[390] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 391) begin
                        n_Body_x[391] = c_Body_x[390];
                        n_Body_y[391] = c_Body_y[390];
                    end else begin
                        n_Body_x[391] = c_Body_x[c_Size-1];
                        n_Body_y[391] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 392) begin
                        n_Body_x[392] = c_Body_x[391];
                        n_Body_y[392] = c_Body_y[391];
                    end else begin
                        n_Body_x[392] = c_Body_x[c_Size-1];
                        n_Body_y[392] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 393) begin
                        n_Body_x[393] = c_Body_x[392];
                        n_Body_y[393] = c_Body_y[392];
                    end else begin
                        n_Body_x[393] = c_Body_x[c_Size-1];
                        n_Body_y[393] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 394) begin
                        n_Body_x[394] = c_Body_x[393];
                        n_Body_y[394] = c_Body_y[393];
                    end else begin
                        n_Body_x[394] = c_Body_x[c_Size-1];
                        n_Body_y[394] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 395) begin
                        n_Body_x[395] = c_Body_x[394];
                        n_Body_y[395] = c_Body_y[394];
                    end else begin
                        n_Body_x[395] = c_Body_x[c_Size-1];
                        n_Body_y[395] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 396) begin
                        n_Body_x[396] = c_Body_x[395];
                        n_Body_y[396] = c_Body_y[395];
                    end else begin
                        n_Body_x[396] = c_Body_x[c_Size-1];
                        n_Body_y[396] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 397) begin
                        n_Body_x[397] = c_Body_x[396];
                        n_Body_y[397] = c_Body_y[396];
                    end else begin
                        n_Body_x[397] = c_Body_x[c_Size-1];
                        n_Body_y[397] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 398) begin
                        n_Body_x[398] = c_Body_x[397];
                        n_Body_y[398] = c_Body_y[397];
                    end else begin
                        n_Body_x[398] = c_Body_x[c_Size-1];
                        n_Body_y[398] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 399) begin
                        n_Body_x[399] = c_Body_x[398];
                        n_Body_y[399] = c_Body_y[398];
                    end else begin
                        n_Body_x[399] = c_Body_x[c_Size-1];
                        n_Body_y[399] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 400) begin
                        n_Body_x[400] = c_Body_x[399];
                        n_Body_y[400] = c_Body_y[399];
                    end else begin
                        n_Body_x[400] = c_Body_x[c_Size-1];
                        n_Body_y[400] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 401) begin
                        n_Body_x[401] = c_Body_x[400];
                        n_Body_y[401] = c_Body_y[400];
                    end else begin
                        n_Body_x[401] = c_Body_x[c_Size-1];
                        n_Body_y[401] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 402) begin
                        n_Body_x[402] = c_Body_x[401];
                        n_Body_y[402] = c_Body_y[401];
                    end else begin
                        n_Body_x[402] = c_Body_x[c_Size-1];
                        n_Body_y[402] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 403) begin
                        n_Body_x[403] = c_Body_x[402];
                        n_Body_y[403] = c_Body_y[402];
                    end else begin
                        n_Body_x[403] = c_Body_x[c_Size-1];
                        n_Body_y[403] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 404) begin
                        n_Body_x[404] = c_Body_x[403];
                        n_Body_y[404] = c_Body_y[403];
                    end else begin
                        n_Body_x[404] = c_Body_x[c_Size-1];
                        n_Body_y[404] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 405) begin
                        n_Body_x[405] = c_Body_x[404];
                        n_Body_y[405] = c_Body_y[404];
                    end else begin
                        n_Body_x[405] = c_Body_x[c_Size-1];
                        n_Body_y[405] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 406) begin
                        n_Body_x[406] = c_Body_x[405];
                        n_Body_y[406] = c_Body_y[405];
                    end else begin
                        n_Body_x[406] = c_Body_x[c_Size-1];
                        n_Body_y[406] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 407) begin
                        n_Body_x[407] = c_Body_x[406];
                        n_Body_y[407] = c_Body_y[406];
                    end else begin
                        n_Body_x[407] = c_Body_x[c_Size-1];
                        n_Body_y[407] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 408) begin
                        n_Body_x[408] = c_Body_x[407];
                        n_Body_y[408] = c_Body_y[407];
                    end else begin
                        n_Body_x[408] = c_Body_x[c_Size-1];
                        n_Body_y[408] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 409) begin
                        n_Body_x[409] = c_Body_x[408];
                        n_Body_y[409] = c_Body_y[408];
                    end else begin
                        n_Body_x[409] = c_Body_x[c_Size-1];
                        n_Body_y[409] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 410) begin
                        n_Body_x[410] = c_Body_x[409];
                        n_Body_y[410] = c_Body_y[409];
                    end else begin
                        n_Body_x[410] = c_Body_x[c_Size-1];
                        n_Body_y[410] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 411) begin
                        n_Body_x[411] = c_Body_x[410];
                        n_Body_y[411] = c_Body_y[410];
                    end else begin
                        n_Body_x[411] = c_Body_x[c_Size-1];
                        n_Body_y[411] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 412) begin
                        n_Body_x[412] = c_Body_x[411];
                        n_Body_y[412] = c_Body_y[411];
                    end else begin
                        n_Body_x[412] = c_Body_x[c_Size-1];
                        n_Body_y[412] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 413) begin
                        n_Body_x[413] = c_Body_x[412];
                        n_Body_y[413] = c_Body_y[412];
                    end else begin
                        n_Body_x[413] = c_Body_x[c_Size-1];
                        n_Body_y[413] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 414) begin
                        n_Body_x[414] = c_Body_x[413];
                        n_Body_y[414] = c_Body_y[413];
                    end else begin
                        n_Body_x[414] = c_Body_x[c_Size-1];
                        n_Body_y[414] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 415) begin
                        n_Body_x[415] = c_Body_x[414];
                        n_Body_y[415] = c_Body_y[414];
                    end else begin
                        n_Body_x[415] = c_Body_x[c_Size-1];
                        n_Body_y[415] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 416) begin
                        n_Body_x[416] = c_Body_x[415];
                        n_Body_y[416] = c_Body_y[415];
                    end else begin
                        n_Body_x[416] = c_Body_x[c_Size-1];
                        n_Body_y[416] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 417) begin
                        n_Body_x[417] = c_Body_x[416];
                        n_Body_y[417] = c_Body_y[416];
                    end else begin
                        n_Body_x[417] = c_Body_x[c_Size-1];
                        n_Body_y[417] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 418) begin
                        n_Body_x[418] = c_Body_x[417];
                        n_Body_y[418] = c_Body_y[417];
                    end else begin
                        n_Body_x[418] = c_Body_x[c_Size-1];
                        n_Body_y[418] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 419) begin
                        n_Body_x[419] = c_Body_x[418];
                        n_Body_y[419] = c_Body_y[418];
                    end else begin
                        n_Body_x[419] = c_Body_x[c_Size-1];
                        n_Body_y[419] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 420) begin
                        n_Body_x[420] = c_Body_x[419];
                        n_Body_y[420] = c_Body_y[419];
                    end else begin
                        n_Body_x[420] = c_Body_x[c_Size-1];
                        n_Body_y[420] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 421) begin
                        n_Body_x[421] = c_Body_x[420];
                        n_Body_y[421] = c_Body_y[420];
                    end else begin
                        n_Body_x[421] = c_Body_x[c_Size-1];
                        n_Body_y[421] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 422) begin
                        n_Body_x[422] = c_Body_x[421];
                        n_Body_y[422] = c_Body_y[421];
                    end else begin
                        n_Body_x[422] = c_Body_x[c_Size-1];
                        n_Body_y[422] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 423) begin
                        n_Body_x[423] = c_Body_x[422];
                        n_Body_y[423] = c_Body_y[422];
                    end else begin
                        n_Body_x[423] = c_Body_x[c_Size-1];
                        n_Body_y[423] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 424) begin
                        n_Body_x[424] = c_Body_x[423];
                        n_Body_y[424] = c_Body_y[423];
                    end else begin
                        n_Body_x[424] = c_Body_x[c_Size-1];
                        n_Body_y[424] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 425) begin
                        n_Body_x[425] = c_Body_x[424];
                        n_Body_y[425] = c_Body_y[424];
                    end else begin
                        n_Body_x[425] = c_Body_x[c_Size-1];
                        n_Body_y[425] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 426) begin
                        n_Body_x[426] = c_Body_x[425];
                        n_Body_y[426] = c_Body_y[425];
                    end else begin
                        n_Body_x[426] = c_Body_x[c_Size-1];
                        n_Body_y[426] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 427) begin
                        n_Body_x[427] = c_Body_x[426];
                        n_Body_y[427] = c_Body_y[426];
                    end else begin
                        n_Body_x[427] = c_Body_x[c_Size-1];
                        n_Body_y[427] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 428) begin
                        n_Body_x[428] = c_Body_x[427];
                        n_Body_y[428] = c_Body_y[427];
                    end else begin
                        n_Body_x[428] = c_Body_x[c_Size-1];
                        n_Body_y[428] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 429) begin
                        n_Body_x[429] = c_Body_x[428];
                        n_Body_y[429] = c_Body_y[428];
                    end else begin
                        n_Body_x[429] = c_Body_x[c_Size-1];
                        n_Body_y[429] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 430) begin
                        n_Body_x[430] = c_Body_x[429];
                        n_Body_y[430] = c_Body_y[429];
                    end else begin
                        n_Body_x[430] = c_Body_x[c_Size-1];
                        n_Body_y[430] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 431) begin
                        n_Body_x[431] = c_Body_x[430];
                        n_Body_y[431] = c_Body_y[430];
                    end else begin
                        n_Body_x[431] = c_Body_x[c_Size-1];
                        n_Body_y[431] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 432) begin
                        n_Body_x[432] = c_Body_x[431];
                        n_Body_y[432] = c_Body_y[431];
                    end else begin
                        n_Body_x[432] = c_Body_x[c_Size-1];
                        n_Body_y[432] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 433) begin
                        n_Body_x[433] = c_Body_x[432];
                        n_Body_y[433] = c_Body_y[432];
                    end else begin
                        n_Body_x[433] = c_Body_x[c_Size-1];
                        n_Body_y[433] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 434) begin
                        n_Body_x[434] = c_Body_x[433];
                        n_Body_y[434] = c_Body_y[433];
                    end else begin
                        n_Body_x[434] = c_Body_x[c_Size-1];
                        n_Body_y[434] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 435) begin
                        n_Body_x[435] = c_Body_x[434];
                        n_Body_y[435] = c_Body_y[434];
                    end else begin
                        n_Body_x[435] = c_Body_x[c_Size-1];
                        n_Body_y[435] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 436) begin
                        n_Body_x[436] = c_Body_x[435];
                        n_Body_y[436] = c_Body_y[435];
                    end else begin
                        n_Body_x[436] = c_Body_x[c_Size-1];
                        n_Body_y[436] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 437) begin
                        n_Body_x[437] = c_Body_x[436];
                        n_Body_y[437] = c_Body_y[436];
                    end else begin
                        n_Body_x[437] = c_Body_x[c_Size-1];
                        n_Body_y[437] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 438) begin
                        n_Body_x[438] = c_Body_x[437];
                        n_Body_y[438] = c_Body_y[437];
                    end else begin
                        n_Body_x[438] = c_Body_x[c_Size-1];
                        n_Body_y[438] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 439) begin
                        n_Body_x[439] = c_Body_x[438];
                        n_Body_y[439] = c_Body_y[438];
                    end else begin
                        n_Body_x[439] = c_Body_x[c_Size-1];
                        n_Body_y[439] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 440) begin
                        n_Body_x[440] = c_Body_x[439];
                        n_Body_y[440] = c_Body_y[439];
                    end else begin
                        n_Body_x[440] = c_Body_x[c_Size-1];
                        n_Body_y[440] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 441) begin
                        n_Body_x[441] = c_Body_x[440];
                        n_Body_y[441] = c_Body_y[440];
                    end else begin
                        n_Body_x[441] = c_Body_x[c_Size-1];
                        n_Body_y[441] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 442) begin
                        n_Body_x[442] = c_Body_x[441];
                        n_Body_y[442] = c_Body_y[441];
                    end else begin
                        n_Body_x[442] = c_Body_x[c_Size-1];
                        n_Body_y[442] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 443) begin
                        n_Body_x[443] = c_Body_x[442];
                        n_Body_y[443] = c_Body_y[442];
                    end else begin
                        n_Body_x[443] = c_Body_x[c_Size-1];
                        n_Body_y[443] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 444) begin
                        n_Body_x[444] = c_Body_x[443];
                        n_Body_y[444] = c_Body_y[443];
                    end else begin
                        n_Body_x[444] = c_Body_x[c_Size-1];
                        n_Body_y[444] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 445) begin
                        n_Body_x[445] = c_Body_x[444];
                        n_Body_y[445] = c_Body_y[444];
                    end else begin
                        n_Body_x[445] = c_Body_x[c_Size-1];
                        n_Body_y[445] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 446) begin
                        n_Body_x[446] = c_Body_x[445];
                        n_Body_y[446] = c_Body_y[445];
                    end else begin
                        n_Body_x[446] = c_Body_x[c_Size-1];
                        n_Body_y[446] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 447) begin
                        n_Body_x[447] = c_Body_x[446];
                        n_Body_y[447] = c_Body_y[446];
                    end else begin
                        n_Body_x[447] = c_Body_x[c_Size-1];
                        n_Body_y[447] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 448) begin
                        n_Body_x[448] = c_Body_x[447];
                        n_Body_y[448] = c_Body_y[447];
                    end else begin
                        n_Body_x[448] = c_Body_x[c_Size-1];
                        n_Body_y[448] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 449) begin
                        n_Body_x[449] = c_Body_x[448];
                        n_Body_y[449] = c_Body_y[448];
                    end else begin
                        n_Body_x[449] = c_Body_x[c_Size-1];
                        n_Body_y[449] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 450) begin
                        n_Body_x[450] = c_Body_x[449];
                        n_Body_y[450] = c_Body_y[449];
                    end else begin
                        n_Body_x[450] = c_Body_x[c_Size-1];
                        n_Body_y[450] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 451) begin
                        n_Body_x[451] = c_Body_x[450];
                        n_Body_y[451] = c_Body_y[450];
                    end else begin
                        n_Body_x[451] = c_Body_x[c_Size-1];
                        n_Body_y[451] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 452) begin
                        n_Body_x[452] = c_Body_x[451];
                        n_Body_y[452] = c_Body_y[451];
                    end else begin
                        n_Body_x[452] = c_Body_x[c_Size-1];
                        n_Body_y[452] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 453) begin
                        n_Body_x[453] = c_Body_x[452];
                        n_Body_y[453] = c_Body_y[452];
                    end else begin
                        n_Body_x[453] = c_Body_x[c_Size-1];
                        n_Body_y[453] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 454) begin
                        n_Body_x[454] = c_Body_x[453];
                        n_Body_y[454] = c_Body_y[453];
                    end else begin
                        n_Body_x[454] = c_Body_x[c_Size-1];
                        n_Body_y[454] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 455) begin
                        n_Body_x[455] = c_Body_x[454];
                        n_Body_y[455] = c_Body_y[454];
                    end else begin
                        n_Body_x[455] = c_Body_x[c_Size-1];
                        n_Body_y[455] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 456) begin
                        n_Body_x[456] = c_Body_x[455];
                        n_Body_y[456] = c_Body_y[455];
                    end else begin
                        n_Body_x[456] = c_Body_x[c_Size-1];
                        n_Body_y[456] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 457) begin
                        n_Body_x[457] = c_Body_x[456];
                        n_Body_y[457] = c_Body_y[456];
                    end else begin
                        n_Body_x[457] = c_Body_x[c_Size-1];
                        n_Body_y[457] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 458) begin
                        n_Body_x[458] = c_Body_x[457];
                        n_Body_y[458] = c_Body_y[457];
                    end else begin
                        n_Body_x[458] = c_Body_x[c_Size-1];
                        n_Body_y[458] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 459) begin
                        n_Body_x[459] = c_Body_x[458];
                        n_Body_y[459] = c_Body_y[458];
                    end else begin
                        n_Body_x[459] = c_Body_x[c_Size-1];
                        n_Body_y[459] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 460) begin
                        n_Body_x[460] = c_Body_x[459];
                        n_Body_y[460] = c_Body_y[459];
                    end else begin
                        n_Body_x[460] = c_Body_x[c_Size-1];
                        n_Body_y[460] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 461) begin
                        n_Body_x[461] = c_Body_x[460];
                        n_Body_y[461] = c_Body_y[460];
                    end else begin
                        n_Body_x[461] = c_Body_x[c_Size-1];
                        n_Body_y[461] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 462) begin
                        n_Body_x[462] = c_Body_x[461];
                        n_Body_y[462] = c_Body_y[461];
                    end else begin
                        n_Body_x[462] = c_Body_x[c_Size-1];
                        n_Body_y[462] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 463) begin
                        n_Body_x[463] = c_Body_x[462];
                        n_Body_y[463] = c_Body_y[462];
                    end else begin
                        n_Body_x[463] = c_Body_x[c_Size-1];
                        n_Body_y[463] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 464) begin
                        n_Body_x[464] = c_Body_x[463];
                        n_Body_y[464] = c_Body_y[463];
                    end else begin
                        n_Body_x[464] = c_Body_x[c_Size-1];
                        n_Body_y[464] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 465) begin
                        n_Body_x[465] = c_Body_x[464];
                        n_Body_y[465] = c_Body_y[464];
                    end else begin
                        n_Body_x[465] = c_Body_x[c_Size-1];
                        n_Body_y[465] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 466) begin
                        n_Body_x[466] = c_Body_x[465];
                        n_Body_y[466] = c_Body_y[465];
                    end else begin
                        n_Body_x[466] = c_Body_x[c_Size-1];
                        n_Body_y[466] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 467) begin
                        n_Body_x[467] = c_Body_x[466];
                        n_Body_y[467] = c_Body_y[466];
                    end else begin
                        n_Body_x[467] = c_Body_x[c_Size-1];
                        n_Body_y[467] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 468) begin
                        n_Body_x[468] = c_Body_x[467];
                        n_Body_y[468] = c_Body_y[467];
                    end else begin
                        n_Body_x[468] = c_Body_x[c_Size-1];
                        n_Body_y[468] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 469) begin
                        n_Body_x[469] = c_Body_x[468];
                        n_Body_y[469] = c_Body_y[468];
                    end else begin
                        n_Body_x[469] = c_Body_x[c_Size-1];
                        n_Body_y[469] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 470) begin
                        n_Body_x[470] = c_Body_x[469];
                        n_Body_y[470] = c_Body_y[469];
                    end else begin
                        n_Body_x[470] = c_Body_x[c_Size-1];
                        n_Body_y[470] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 471) begin
                        n_Body_x[471] = c_Body_x[470];
                        n_Body_y[471] = c_Body_y[470];
                    end else begin
                        n_Body_x[471] = c_Body_x[c_Size-1];
                        n_Body_y[471] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 472) begin
                        n_Body_x[472] = c_Body_x[471];
                        n_Body_y[472] = c_Body_y[471];
                    end else begin
                        n_Body_x[472] = c_Body_x[c_Size-1];
                        n_Body_y[472] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 473) begin
                        n_Body_x[473] = c_Body_x[472];
                        n_Body_y[473] = c_Body_y[472];
                    end else begin
                        n_Body_x[473] = c_Body_x[c_Size-1];
                        n_Body_y[473] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 474) begin
                        n_Body_x[474] = c_Body_x[473];
                        n_Body_y[474] = c_Body_y[473];
                    end else begin
                        n_Body_x[474] = c_Body_x[c_Size-1];
                        n_Body_y[474] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 475) begin
                        n_Body_x[475] = c_Body_x[474];
                        n_Body_y[475] = c_Body_y[474];
                    end else begin
                        n_Body_x[475] = c_Body_x[c_Size-1];
                        n_Body_y[475] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 476) begin
                        n_Body_x[476] = c_Body_x[475];
                        n_Body_y[476] = c_Body_y[475];
                    end else begin
                        n_Body_x[476] = c_Body_x[c_Size-1];
                        n_Body_y[476] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 477) begin
                        n_Body_x[477] = c_Body_x[476];
                        n_Body_y[477] = c_Body_y[476];
                    end else begin
                        n_Body_x[477] = c_Body_x[c_Size-1];
                        n_Body_y[477] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 478) begin
                        n_Body_x[478] = c_Body_x[477];
                        n_Body_y[478] = c_Body_y[477];
                    end else begin
                        n_Body_x[478] = c_Body_x[c_Size-1];
                        n_Body_y[478] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 479) begin
                        n_Body_x[479] = c_Body_x[478];
                        n_Body_y[479] = c_Body_y[478];
                    end else begin
                        n_Body_x[479] = c_Body_x[c_Size-1];
                        n_Body_y[479] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 480) begin
                        n_Body_x[480] = c_Body_x[479];
                        n_Body_y[480] = c_Body_y[479];
                    end else begin
                        n_Body_x[480] = c_Body_x[c_Size-1];
                        n_Body_y[480] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 481) begin
                        n_Body_x[481] = c_Body_x[480];
                        n_Body_y[481] = c_Body_y[480];
                    end else begin
                        n_Body_x[481] = c_Body_x[c_Size-1];
                        n_Body_y[481] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 482) begin
                        n_Body_x[482] = c_Body_x[481];
                        n_Body_y[482] = c_Body_y[481];
                    end else begin
                        n_Body_x[482] = c_Body_x[c_Size-1];
                        n_Body_y[482] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 483) begin
                        n_Body_x[483] = c_Body_x[482];
                        n_Body_y[483] = c_Body_y[482];
                    end else begin
                        n_Body_x[483] = c_Body_x[c_Size-1];
                        n_Body_y[483] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 484) begin
                        n_Body_x[484] = c_Body_x[483];
                        n_Body_y[484] = c_Body_y[483];
                    end else begin
                        n_Body_x[484] = c_Body_x[c_Size-1];
                        n_Body_y[484] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 485) begin
                        n_Body_x[485] = c_Body_x[484];
                        n_Body_y[485] = c_Body_y[484];
                    end else begin
                        n_Body_x[485] = c_Body_x[c_Size-1];
                        n_Body_y[485] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 486) begin
                        n_Body_x[486] = c_Body_x[485];
                        n_Body_y[486] = c_Body_y[485];
                    end else begin
                        n_Body_x[486] = c_Body_x[c_Size-1];
                        n_Body_y[486] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 487) begin
                        n_Body_x[487] = c_Body_x[486];
                        n_Body_y[487] = c_Body_y[486];
                    end else begin
                        n_Body_x[487] = c_Body_x[c_Size-1];
                        n_Body_y[487] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 488) begin
                        n_Body_x[488] = c_Body_x[487];
                        n_Body_y[488] = c_Body_y[487];
                    end else begin
                        n_Body_x[488] = c_Body_x[c_Size-1];
                        n_Body_y[488] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 489) begin
                        n_Body_x[489] = c_Body_x[488];
                        n_Body_y[489] = c_Body_y[488];
                    end else begin
                        n_Body_x[489] = c_Body_x[c_Size-1];
                        n_Body_y[489] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 490) begin
                        n_Body_x[490] = c_Body_x[489];
                        n_Body_y[490] = c_Body_y[489];
                    end else begin
                        n_Body_x[490] = c_Body_x[c_Size-1];
                        n_Body_y[490] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 491) begin
                        n_Body_x[491] = c_Body_x[490];
                        n_Body_y[491] = c_Body_y[490];
                    end else begin
                        n_Body_x[491] = c_Body_x[c_Size-1];
                        n_Body_y[491] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 492) begin
                        n_Body_x[492] = c_Body_x[491];
                        n_Body_y[492] = c_Body_y[491];
                    end else begin
                        n_Body_x[492] = c_Body_x[c_Size-1];
                        n_Body_y[492] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 493) begin
                        n_Body_x[493] = c_Body_x[492];
                        n_Body_y[493] = c_Body_y[492];
                    end else begin
                        n_Body_x[493] = c_Body_x[c_Size-1];
                        n_Body_y[493] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 494) begin
                        n_Body_x[494] = c_Body_x[493];
                        n_Body_y[494] = c_Body_y[493];
                    end else begin
                        n_Body_x[494] = c_Body_x[c_Size-1];
                        n_Body_y[494] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 495) begin
                        n_Body_x[495] = c_Body_x[494];
                        n_Body_y[495] = c_Body_y[494];
                    end else begin
                        n_Body_x[495] = c_Body_x[c_Size-1];
                        n_Body_y[495] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 496) begin
                        n_Body_x[496] = c_Body_x[495];
                        n_Body_y[496] = c_Body_y[495];
                    end else begin
                        n_Body_x[496] = c_Body_x[c_Size-1];
                        n_Body_y[496] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 497) begin
                        n_Body_x[497] = c_Body_x[496];
                        n_Body_y[497] = c_Body_y[496];
                    end else begin
                        n_Body_x[497] = c_Body_x[c_Size-1];
                        n_Body_y[497] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 498) begin
                        n_Body_x[498] = c_Body_x[497];
                        n_Body_y[498] = c_Body_y[497];
                    end else begin
                        n_Body_x[498] = c_Body_x[c_Size-1];
                        n_Body_y[498] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 499) begin
                        n_Body_x[499] = c_Body_x[498];
                        n_Body_y[499] = c_Body_y[498];
                    end else begin
                        n_Body_x[499] = c_Body_x[c_Size-1];
                        n_Body_y[499] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 500) begin
                        n_Body_x[500] = c_Body_x[499];
                        n_Body_y[500] = c_Body_y[499];
                    end else begin
                        n_Body_x[500] = c_Body_x[c_Size-1];
                        n_Body_y[500] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 501) begin
                        n_Body_x[501] = c_Body_x[500];
                        n_Body_y[501] = c_Body_y[500];
                    end else begin
                        n_Body_x[501] = c_Body_x[c_Size-1];
                        n_Body_y[501] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 502) begin
                        n_Body_x[502] = c_Body_x[501];
                        n_Body_y[502] = c_Body_y[501];
                    end else begin
                        n_Body_x[502] = c_Body_x[c_Size-1];
                        n_Body_y[502] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 503) begin
                        n_Body_x[503] = c_Body_x[502];
                        n_Body_y[503] = c_Body_y[502];
                    end else begin
                        n_Body_x[503] = c_Body_x[c_Size-1];
                        n_Body_y[503] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 504) begin
                        n_Body_x[504] = c_Body_x[503];
                        n_Body_y[504] = c_Body_y[503];
                    end else begin
                        n_Body_x[504] = c_Body_x[c_Size-1];
                        n_Body_y[504] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 505) begin
                        n_Body_x[505] = c_Body_x[504];
                        n_Body_y[505] = c_Body_y[504];
                    end else begin
                        n_Body_x[505] = c_Body_x[c_Size-1];
                        n_Body_y[505] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 506) begin
                        n_Body_x[506] = c_Body_x[505];
                        n_Body_y[506] = c_Body_y[505];
                    end else begin
                        n_Body_x[506] = c_Body_x[c_Size-1];
                        n_Body_y[506] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 507) begin
                        n_Body_x[507] = c_Body_x[506];
                        n_Body_y[507] = c_Body_y[506];
                    end else begin
                        n_Body_x[507] = c_Body_x[c_Size-1];
                        n_Body_y[507] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 508) begin
                        n_Body_x[508] = c_Body_x[507];
                        n_Body_y[508] = c_Body_y[507];
                    end else begin
                        n_Body_x[508] = c_Body_x[c_Size-1];
                        n_Body_y[508] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 509) begin
                        n_Body_x[509] = c_Body_x[508];
                        n_Body_y[509] = c_Body_y[508];
                    end else begin
                        n_Body_x[509] = c_Body_x[c_Size-1];
                        n_Body_y[509] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 510) begin
                        n_Body_x[510] = c_Body_x[509];
                        n_Body_y[510] = c_Body_y[509];
                    end else begin
                        n_Body_x[510] = c_Body_x[c_Size-1];
                        n_Body_y[510] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 511) begin
                        n_Body_x[511] = c_Body_x[510];
                        n_Body_y[511] = c_Body_y[510];
                    end else begin
                        n_Body_x[511] = c_Body_x[c_Size-1];
                        n_Body_y[511] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 512) begin
                        n_Body_x[512] = c_Body_x[511];
                        n_Body_y[512] = c_Body_y[511];
                    end else begin
                        n_Body_x[512] = c_Body_x[c_Size-1];
                        n_Body_y[512] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 513) begin
                        n_Body_x[513] = c_Body_x[512];
                        n_Body_y[513] = c_Body_y[512];
                    end else begin
                        n_Body_x[513] = c_Body_x[c_Size-1];
                        n_Body_y[513] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 514) begin
                        n_Body_x[514] = c_Body_x[513];
                        n_Body_y[514] = c_Body_y[513];
                    end else begin
                        n_Body_x[514] = c_Body_x[c_Size-1];
                        n_Body_y[514] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 515) begin
                        n_Body_x[515] = c_Body_x[514];
                        n_Body_y[515] = c_Body_y[514];
                    end else begin
                        n_Body_x[515] = c_Body_x[c_Size-1];
                        n_Body_y[515] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 516) begin
                        n_Body_x[516] = c_Body_x[515];
                        n_Body_y[516] = c_Body_y[515];
                    end else begin
                        n_Body_x[516] = c_Body_x[c_Size-1];
                        n_Body_y[516] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 517) begin
                        n_Body_x[517] = c_Body_x[516];
                        n_Body_y[517] = c_Body_y[516];
                    end else begin
                        n_Body_x[517] = c_Body_x[c_Size-1];
                        n_Body_y[517] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 518) begin
                        n_Body_x[518] = c_Body_x[517];
                        n_Body_y[518] = c_Body_y[517];
                    end else begin
                        n_Body_x[518] = c_Body_x[c_Size-1];
                        n_Body_y[518] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 519) begin
                        n_Body_x[519] = c_Body_x[518];
                        n_Body_y[519] = c_Body_y[518];
                    end else begin
                        n_Body_x[519] = c_Body_x[c_Size-1];
                        n_Body_y[519] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 520) begin
                        n_Body_x[520] = c_Body_x[519];
                        n_Body_y[520] = c_Body_y[519];
                    end else begin
                        n_Body_x[520] = c_Body_x[c_Size-1];
                        n_Body_y[520] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 521) begin
                        n_Body_x[521] = c_Body_x[520];
                        n_Body_y[521] = c_Body_y[520];
                    end else begin
                        n_Body_x[521] = c_Body_x[c_Size-1];
                        n_Body_y[521] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 522) begin
                        n_Body_x[522] = c_Body_x[521];
                        n_Body_y[522] = c_Body_y[521];
                    end else begin
                        n_Body_x[522] = c_Body_x[c_Size-1];
                        n_Body_y[522] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 523) begin
                        n_Body_x[523] = c_Body_x[522];
                        n_Body_y[523] = c_Body_y[522];
                    end else begin
                        n_Body_x[523] = c_Body_x[c_Size-1];
                        n_Body_y[523] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 524) begin
                        n_Body_x[524] = c_Body_x[523];
                        n_Body_y[524] = c_Body_y[523];
                    end else begin
                        n_Body_x[524] = c_Body_x[c_Size-1];
                        n_Body_y[524] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 525) begin
                        n_Body_x[525] = c_Body_x[524];
                        n_Body_y[525] = c_Body_y[524];
                    end else begin
                        n_Body_x[525] = c_Body_x[c_Size-1];
                        n_Body_y[525] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 526) begin
                        n_Body_x[526] = c_Body_x[525];
                        n_Body_y[526] = c_Body_y[525];
                    end else begin
                        n_Body_x[526] = c_Body_x[c_Size-1];
                        n_Body_y[526] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 527) begin
                        n_Body_x[527] = c_Body_x[526];
                        n_Body_y[527] = c_Body_y[526];
                    end else begin
                        n_Body_x[527] = c_Body_x[c_Size-1];
                        n_Body_y[527] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 528) begin
                        n_Body_x[528] = c_Body_x[527];
                        n_Body_y[528] = c_Body_y[527];
                    end else begin
                        n_Body_x[528] = c_Body_x[c_Size-1];
                        n_Body_y[528] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 529) begin
                        n_Body_x[529] = c_Body_x[528];
                        n_Body_y[529] = c_Body_y[528];
                    end else begin
                        n_Body_x[529] = c_Body_x[c_Size-1];
                        n_Body_y[529] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 530) begin
                        n_Body_x[530] = c_Body_x[529];
                        n_Body_y[530] = c_Body_y[529];
                    end else begin
                        n_Body_x[530] = c_Body_x[c_Size-1];
                        n_Body_y[530] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 531) begin
                        n_Body_x[531] = c_Body_x[530];
                        n_Body_y[531] = c_Body_y[530];
                    end else begin
                        n_Body_x[531] = c_Body_x[c_Size-1];
                        n_Body_y[531] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 532) begin
                        n_Body_x[532] = c_Body_x[531];
                        n_Body_y[532] = c_Body_y[531];
                    end else begin
                        n_Body_x[532] = c_Body_x[c_Size-1];
                        n_Body_y[532] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 533) begin
                        n_Body_x[533] = c_Body_x[532];
                        n_Body_y[533] = c_Body_y[532];
                    end else begin
                        n_Body_x[533] = c_Body_x[c_Size-1];
                        n_Body_y[533] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 534) begin
                        n_Body_x[534] = c_Body_x[533];
                        n_Body_y[534] = c_Body_y[533];
                    end else begin
                        n_Body_x[534] = c_Body_x[c_Size-1];
                        n_Body_y[534] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 535) begin
                        n_Body_x[535] = c_Body_x[534];
                        n_Body_y[535] = c_Body_y[534];
                    end else begin
                        n_Body_x[535] = c_Body_x[c_Size-1];
                        n_Body_y[535] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 536) begin
                        n_Body_x[536] = c_Body_x[535];
                        n_Body_y[536] = c_Body_y[535];
                    end else begin
                        n_Body_x[536] = c_Body_x[c_Size-1];
                        n_Body_y[536] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 537) begin
                        n_Body_x[537] = c_Body_x[536];
                        n_Body_y[537] = c_Body_y[536];
                    end else begin
                        n_Body_x[537] = c_Body_x[c_Size-1];
                        n_Body_y[537] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 538) begin
                        n_Body_x[538] = c_Body_x[537];
                        n_Body_y[538] = c_Body_y[537];
                    end else begin
                        n_Body_x[538] = c_Body_x[c_Size-1];
                        n_Body_y[538] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 539) begin
                        n_Body_x[539] = c_Body_x[538];
                        n_Body_y[539] = c_Body_y[538];
                    end else begin
                        n_Body_x[539] = c_Body_x[c_Size-1];
                        n_Body_y[539] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 540) begin
                        n_Body_x[540] = c_Body_x[539];
                        n_Body_y[540] = c_Body_y[539];
                    end else begin
                        n_Body_x[540] = c_Body_x[c_Size-1];
                        n_Body_y[540] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 541) begin
                        n_Body_x[541] = c_Body_x[540];
                        n_Body_y[541] = c_Body_y[540];
                    end else begin
                        n_Body_x[541] = c_Body_x[c_Size-1];
                        n_Body_y[541] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 542) begin
                        n_Body_x[542] = c_Body_x[541];
                        n_Body_y[542] = c_Body_y[541];
                    end else begin
                        n_Body_x[542] = c_Body_x[c_Size-1];
                        n_Body_y[542] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 543) begin
                        n_Body_x[543] = c_Body_x[542];
                        n_Body_y[543] = c_Body_y[542];
                    end else begin
                        n_Body_x[543] = c_Body_x[c_Size-1];
                        n_Body_y[543] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 544) begin
                        n_Body_x[544] = c_Body_x[543];
                        n_Body_y[544] = c_Body_y[543];
                    end else begin
                        n_Body_x[544] = c_Body_x[c_Size-1];
                        n_Body_y[544] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 545) begin
                        n_Body_x[545] = c_Body_x[544];
                        n_Body_y[545] = c_Body_y[544];
                    end else begin
                        n_Body_x[545] = c_Body_x[c_Size-1];
                        n_Body_y[545] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 546) begin
                        n_Body_x[546] = c_Body_x[545];
                        n_Body_y[546] = c_Body_y[545];
                    end else begin
                        n_Body_x[546] = c_Body_x[c_Size-1];
                        n_Body_y[546] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 547) begin
                        n_Body_x[547] = c_Body_x[546];
                        n_Body_y[547] = c_Body_y[546];
                    end else begin
                        n_Body_x[547] = c_Body_x[c_Size-1];
                        n_Body_y[547] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 548) begin
                        n_Body_x[548] = c_Body_x[547];
                        n_Body_y[548] = c_Body_y[547];
                    end else begin
                        n_Body_x[548] = c_Body_x[c_Size-1];
                        n_Body_y[548] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 549) begin
                        n_Body_x[549] = c_Body_x[548];
                        n_Body_y[549] = c_Body_y[548];
                    end else begin
                        n_Body_x[549] = c_Body_x[c_Size-1];
                        n_Body_y[549] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 550) begin
                        n_Body_x[550] = c_Body_x[549];
                        n_Body_y[550] = c_Body_y[549];
                    end else begin
                        n_Body_x[550] = c_Body_x[c_Size-1];
                        n_Body_y[550] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 551) begin
                        n_Body_x[551] = c_Body_x[550];
                        n_Body_y[551] = c_Body_y[550];
                    end else begin
                        n_Body_x[551] = c_Body_x[c_Size-1];
                        n_Body_y[551] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 552) begin
                        n_Body_x[552] = c_Body_x[551];
                        n_Body_y[552] = c_Body_y[551];
                    end else begin
                        n_Body_x[552] = c_Body_x[c_Size-1];
                        n_Body_y[552] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 553) begin
                        n_Body_x[553] = c_Body_x[552];
                        n_Body_y[553] = c_Body_y[552];
                    end else begin
                        n_Body_x[553] = c_Body_x[c_Size-1];
                        n_Body_y[553] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 554) begin
                        n_Body_x[554] = c_Body_x[553];
                        n_Body_y[554] = c_Body_y[553];
                    end else begin
                        n_Body_x[554] = c_Body_x[c_Size-1];
                        n_Body_y[554] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 555) begin
                        n_Body_x[555] = c_Body_x[554];
                        n_Body_y[555] = c_Body_y[554];
                    end else begin
                        n_Body_x[555] = c_Body_x[c_Size-1];
                        n_Body_y[555] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 556) begin
                        n_Body_x[556] = c_Body_x[555];
                        n_Body_y[556] = c_Body_y[555];
                    end else begin
                        n_Body_x[556] = c_Body_x[c_Size-1];
                        n_Body_y[556] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 557) begin
                        n_Body_x[557] = c_Body_x[556];
                        n_Body_y[557] = c_Body_y[556];
                    end else begin
                        n_Body_x[557] = c_Body_x[c_Size-1];
                        n_Body_y[557] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 558) begin
                        n_Body_x[558] = c_Body_x[557];
                        n_Body_y[558] = c_Body_y[557];
                    end else begin
                        n_Body_x[558] = c_Body_x[c_Size-1];
                        n_Body_y[558] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 559) begin
                        n_Body_x[559] = c_Body_x[558];
                        n_Body_y[559] = c_Body_y[558];
                    end else begin
                        n_Body_x[559] = c_Body_x[c_Size-1];
                        n_Body_y[559] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 560) begin
                        n_Body_x[560] = c_Body_x[559];
                        n_Body_y[560] = c_Body_y[559];
                    end else begin
                        n_Body_x[560] = c_Body_x[c_Size-1];
                        n_Body_y[560] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 561) begin
                        n_Body_x[561] = c_Body_x[560];
                        n_Body_y[561] = c_Body_y[560];
                    end else begin
                        n_Body_x[561] = c_Body_x[c_Size-1];
                        n_Body_y[561] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 562) begin
                        n_Body_x[562] = c_Body_x[561];
                        n_Body_y[562] = c_Body_y[561];
                    end else begin
                        n_Body_x[562] = c_Body_x[c_Size-1];
                        n_Body_y[562] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 563) begin
                        n_Body_x[563] = c_Body_x[562];
                        n_Body_y[563] = c_Body_y[562];
                    end else begin
                        n_Body_x[563] = c_Body_x[c_Size-1];
                        n_Body_y[563] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 564) begin
                        n_Body_x[564] = c_Body_x[563];
                        n_Body_y[564] = c_Body_y[563];
                    end else begin
                        n_Body_x[564] = c_Body_x[c_Size-1];
                        n_Body_y[564] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 565) begin
                        n_Body_x[565] = c_Body_x[564];
                        n_Body_y[565] = c_Body_y[564];
                    end else begin
                        n_Body_x[565] = c_Body_x[c_Size-1];
                        n_Body_y[565] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 566) begin
                        n_Body_x[566] = c_Body_x[565];
                        n_Body_y[566] = c_Body_y[565];
                    end else begin
                        n_Body_x[566] = c_Body_x[c_Size-1];
                        n_Body_y[566] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 567) begin
                        n_Body_x[567] = c_Body_x[566];
                        n_Body_y[567] = c_Body_y[566];
                    end else begin
                        n_Body_x[567] = c_Body_x[c_Size-1];
                        n_Body_y[567] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 568) begin
                        n_Body_x[568] = c_Body_x[567];
                        n_Body_y[568] = c_Body_y[567];
                    end else begin
                        n_Body_x[568] = c_Body_x[c_Size-1];
                        n_Body_y[568] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 569) begin
                        n_Body_x[569] = c_Body_x[568];
                        n_Body_y[569] = c_Body_y[568];
                    end else begin
                        n_Body_x[569] = c_Body_x[c_Size-1];
                        n_Body_y[569] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 570) begin
                        n_Body_x[570] = c_Body_x[569];
                        n_Body_y[570] = c_Body_y[569];
                    end else begin
                        n_Body_x[570] = c_Body_x[c_Size-1];
                        n_Body_y[570] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 571) begin
                        n_Body_x[571] = c_Body_x[570];
                        n_Body_y[571] = c_Body_y[570];
                    end else begin
                        n_Body_x[571] = c_Body_x[c_Size-1];
                        n_Body_y[571] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 572) begin
                        n_Body_x[572] = c_Body_x[571];
                        n_Body_y[572] = c_Body_y[571];
                    end else begin
                        n_Body_x[572] = c_Body_x[c_Size-1];
                        n_Body_y[572] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 573) begin
                        n_Body_x[573] = c_Body_x[572];
                        n_Body_y[573] = c_Body_y[572];
                    end else begin
                        n_Body_x[573] = c_Body_x[c_Size-1];
                        n_Body_y[573] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 574) begin
                        n_Body_x[574] = c_Body_x[573];
                        n_Body_y[574] = c_Body_y[573];
                    end else begin
                        n_Body_x[574] = c_Body_x[c_Size-1];
                        n_Body_y[574] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 575) begin
                        n_Body_x[575] = c_Body_x[574];
                        n_Body_y[575] = c_Body_y[574];
                    end else begin
                        n_Body_x[575] = c_Body_x[c_Size-1];
                        n_Body_y[575] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 576) begin
                        n_Body_x[576] = c_Body_x[575];
                        n_Body_y[576] = c_Body_y[575];
                    end else begin
                        n_Body_x[576] = c_Body_x[c_Size-1];
                        n_Body_y[576] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 577) begin
                        n_Body_x[577] = c_Body_x[576];
                        n_Body_y[577] = c_Body_y[576];
                    end else begin
                        n_Body_x[577] = c_Body_x[c_Size-1];
                        n_Body_y[577] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 578) begin
                        n_Body_x[578] = c_Body_x[577];
                        n_Body_y[578] = c_Body_y[577];
                    end else begin
                        n_Body_x[578] = c_Body_x[c_Size-1];
                        n_Body_y[578] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 579) begin
                        n_Body_x[579] = c_Body_x[578];
                        n_Body_y[579] = c_Body_y[578];
                    end else begin
                        n_Body_x[579] = c_Body_x[c_Size-1];
                        n_Body_y[579] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 580) begin
                        n_Body_x[580] = c_Body_x[579];
                        n_Body_y[580] = c_Body_y[579];
                    end else begin
                        n_Body_x[580] = c_Body_x[c_Size-1];
                        n_Body_y[580] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 581) begin
                        n_Body_x[581] = c_Body_x[580];
                        n_Body_y[581] = c_Body_y[580];
                    end else begin
                        n_Body_x[581] = c_Body_x[c_Size-1];
                        n_Body_y[581] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 582) begin
                        n_Body_x[582] = c_Body_x[581];
                        n_Body_y[582] = c_Body_y[581];
                    end else begin
                        n_Body_x[582] = c_Body_x[c_Size-1];
                        n_Body_y[582] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 583) begin
                        n_Body_x[583] = c_Body_x[582];
                        n_Body_y[583] = c_Body_y[582];
                    end else begin
                        n_Body_x[583] = c_Body_x[c_Size-1];
                        n_Body_y[583] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 584) begin
                        n_Body_x[584] = c_Body_x[583];
                        n_Body_y[584] = c_Body_y[583];
                    end else begin
                        n_Body_x[584] = c_Body_x[c_Size-1];
                        n_Body_y[584] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 585) begin
                        n_Body_x[585] = c_Body_x[584];
                        n_Body_y[585] = c_Body_y[584];
                    end else begin
                        n_Body_x[585] = c_Body_x[c_Size-1];
                        n_Body_y[585] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 586) begin
                        n_Body_x[586] = c_Body_x[585];
                        n_Body_y[586] = c_Body_y[585];
                    end else begin
                        n_Body_x[586] = c_Body_x[c_Size-1];
                        n_Body_y[586] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 587) begin
                        n_Body_x[587] = c_Body_x[586];
                        n_Body_y[587] = c_Body_y[586];
                    end else begin
                        n_Body_x[587] = c_Body_x[c_Size-1];
                        n_Body_y[587] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 588) begin
                        n_Body_x[588] = c_Body_x[587];
                        n_Body_y[588] = c_Body_y[587];
                    end else begin
                        n_Body_x[588] = c_Body_x[c_Size-1];
                        n_Body_y[588] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 589) begin
                        n_Body_x[589] = c_Body_x[588];
                        n_Body_y[589] = c_Body_y[588];
                    end else begin
                        n_Body_x[589] = c_Body_x[c_Size-1];
                        n_Body_y[589] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 590) begin
                        n_Body_x[590] = c_Body_x[589];
                        n_Body_y[590] = c_Body_y[589];
                    end else begin
                        n_Body_x[590] = c_Body_x[c_Size-1];
                        n_Body_y[590] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 591) begin
                        n_Body_x[591] = c_Body_x[590];
                        n_Body_y[591] = c_Body_y[590];
                    end else begin
                        n_Body_x[591] = c_Body_x[c_Size-1];
                        n_Body_y[591] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 592) begin
                        n_Body_x[592] = c_Body_x[591];
                        n_Body_y[592] = c_Body_y[591];
                    end else begin
                        n_Body_x[592] = c_Body_x[c_Size-1];
                        n_Body_y[592] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 593) begin
                        n_Body_x[593] = c_Body_x[592];
                        n_Body_y[593] = c_Body_y[592];
                    end else begin
                        n_Body_x[593] = c_Body_x[c_Size-1];
                        n_Body_y[593] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 594) begin
                        n_Body_x[594] = c_Body_x[593];
                        n_Body_y[594] = c_Body_y[593];
                    end else begin
                        n_Body_x[594] = c_Body_x[c_Size-1];
                        n_Body_y[594] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 595) begin
                        n_Body_x[595] = c_Body_x[594];
                        n_Body_y[595] = c_Body_y[594];
                    end else begin
                        n_Body_x[595] = c_Body_x[c_Size-1];
                        n_Body_y[595] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 596) begin
                        n_Body_x[596] = c_Body_x[595];
                        n_Body_y[596] = c_Body_y[595];
                    end else begin
                        n_Body_x[596] = c_Body_x[c_Size-1];
                        n_Body_y[596] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 597) begin
                        n_Body_x[597] = c_Body_x[596];
                        n_Body_y[597] = c_Body_y[596];
                    end else begin
                        n_Body_x[597] = c_Body_x[c_Size-1];
                        n_Body_y[597] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 598) begin
                        n_Body_x[598] = c_Body_x[597];
                        n_Body_y[598] = c_Body_y[597];
                    end else begin
                        n_Body_x[598] = c_Body_x[c_Size-1];
                        n_Body_y[598] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 599) begin
                        n_Body_x[599] = c_Body_x[598];
                        n_Body_y[599] = c_Body_y[598];
                    end else begin
                        n_Body_x[599] = c_Body_x[c_Size-1];
                        n_Body_y[599] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 600) begin
                        n_Body_x[600] = c_Body_x[599];
                        n_Body_y[600] = c_Body_y[599];
                    end else begin
                        n_Body_x[600] = c_Body_x[c_Size-1];
                        n_Body_y[600] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 601) begin
                        n_Body_x[601] = c_Body_x[600];
                        n_Body_y[601] = c_Body_y[600];
                    end else begin
                        n_Body_x[601] = c_Body_x[c_Size-1];
                        n_Body_y[601] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 602) begin
                        n_Body_x[602] = c_Body_x[601];
                        n_Body_y[602] = c_Body_y[601];
                    end else begin
                        n_Body_x[602] = c_Body_x[c_Size-1];
                        n_Body_y[602] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 603) begin
                        n_Body_x[603] = c_Body_x[602];
                        n_Body_y[603] = c_Body_y[602];
                    end else begin
                        n_Body_x[603] = c_Body_x[c_Size-1];
                        n_Body_y[603] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 604) begin
                        n_Body_x[604] = c_Body_x[603];
                        n_Body_y[604] = c_Body_y[603];
                    end else begin
                        n_Body_x[604] = c_Body_x[c_Size-1];
                        n_Body_y[604] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 605) begin
                        n_Body_x[605] = c_Body_x[604];
                        n_Body_y[605] = c_Body_y[604];
                    end else begin
                        n_Body_x[605] = c_Body_x[c_Size-1];
                        n_Body_y[605] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 606) begin
                        n_Body_x[606] = c_Body_x[605];
                        n_Body_y[606] = c_Body_y[605];
                    end else begin
                        n_Body_x[606] = c_Body_x[c_Size-1];
                        n_Body_y[606] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 607) begin
                        n_Body_x[607] = c_Body_x[606];
                        n_Body_y[607] = c_Body_y[606];
                    end else begin
                        n_Body_x[607] = c_Body_x[c_Size-1];
                        n_Body_y[607] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 608) begin
                        n_Body_x[608] = c_Body_x[607];
                        n_Body_y[608] = c_Body_y[607];
                    end else begin
                        n_Body_x[608] = c_Body_x[c_Size-1];
                        n_Body_y[608] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 609) begin
                        n_Body_x[609] = c_Body_x[608];
                        n_Body_y[609] = c_Body_y[608];
                    end else begin
                        n_Body_x[609] = c_Body_x[c_Size-1];
                        n_Body_y[609] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 610) begin
                        n_Body_x[610] = c_Body_x[609];
                        n_Body_y[610] = c_Body_y[609];
                    end else begin
                        n_Body_x[610] = c_Body_x[c_Size-1];
                        n_Body_y[610] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 611) begin
                        n_Body_x[611] = c_Body_x[610];
                        n_Body_y[611] = c_Body_y[610];
                    end else begin
                        n_Body_x[611] = c_Body_x[c_Size-1];
                        n_Body_y[611] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 612) begin
                        n_Body_x[612] = c_Body_x[611];
                        n_Body_y[612] = c_Body_y[611];
                    end else begin
                        n_Body_x[612] = c_Body_x[c_Size-1];
                        n_Body_y[612] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 613) begin
                        n_Body_x[613] = c_Body_x[612];
                        n_Body_y[613] = c_Body_y[612];
                    end else begin
                        n_Body_x[613] = c_Body_x[c_Size-1];
                        n_Body_y[613] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 614) begin
                        n_Body_x[614] = c_Body_x[613];
                        n_Body_y[614] = c_Body_y[613];
                    end else begin
                        n_Body_x[614] = c_Body_x[c_Size-1];
                        n_Body_y[614] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 615) begin
                        n_Body_x[615] = c_Body_x[614];
                        n_Body_y[615] = c_Body_y[614];
                    end else begin
                        n_Body_x[615] = c_Body_x[c_Size-1];
                        n_Body_y[615] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 616) begin
                        n_Body_x[616] = c_Body_x[615];
                        n_Body_y[616] = c_Body_y[615];
                    end else begin
                        n_Body_x[616] = c_Body_x[c_Size-1];
                        n_Body_y[616] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 617) begin
                        n_Body_x[617] = c_Body_x[616];
                        n_Body_y[617] = c_Body_y[616];
                    end else begin
                        n_Body_x[617] = c_Body_x[c_Size-1];
                        n_Body_y[617] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 618) begin
                        n_Body_x[618] = c_Body_x[617];
                        n_Body_y[618] = c_Body_y[617];
                    end else begin
                        n_Body_x[618] = c_Body_x[c_Size-1];
                        n_Body_y[618] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 619) begin
                        n_Body_x[619] = c_Body_x[618];
                        n_Body_y[619] = c_Body_y[618];
                    end else begin
                        n_Body_x[619] = c_Body_x[c_Size-1];
                        n_Body_y[619] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 620) begin
                        n_Body_x[620] = c_Body_x[619];
                        n_Body_y[620] = c_Body_y[619];
                    end else begin
                        n_Body_x[620] = c_Body_x[c_Size-1];
                        n_Body_y[620] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 621) begin
                        n_Body_x[621] = c_Body_x[620];
                        n_Body_y[621] = c_Body_y[620];
                    end else begin
                        n_Body_x[621] = c_Body_x[c_Size-1];
                        n_Body_y[621] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 622) begin
                        n_Body_x[622] = c_Body_x[621];
                        n_Body_y[622] = c_Body_y[621];
                    end else begin
                        n_Body_x[622] = c_Body_x[c_Size-1];
                        n_Body_y[622] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 623) begin
                        n_Body_x[623] = c_Body_x[622];
                        n_Body_y[623] = c_Body_y[622];
                    end else begin
                        n_Body_x[623] = c_Body_x[c_Size-1];
                        n_Body_y[623] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 624) begin
                        n_Body_x[624] = c_Body_x[623];
                        n_Body_y[624] = c_Body_y[623];
                    end else begin
                        n_Body_x[624] = c_Body_x[c_Size-1];
                        n_Body_y[624] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 625) begin
                        n_Body_x[625] = c_Body_x[624];
                        n_Body_y[625] = c_Body_y[624];
                    end else begin
                        n_Body_x[625] = c_Body_x[c_Size-1];
                        n_Body_y[625] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 626) begin
                        n_Body_x[626] = c_Body_x[625];
                        n_Body_y[626] = c_Body_y[625];
                    end else begin
                        n_Body_x[626] = c_Body_x[c_Size-1];
                        n_Body_y[626] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 627) begin
                        n_Body_x[627] = c_Body_x[626];
                        n_Body_y[627] = c_Body_y[626];
                    end else begin
                        n_Body_x[627] = c_Body_x[c_Size-1];
                        n_Body_y[627] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 628) begin
                        n_Body_x[628] = c_Body_x[627];
                        n_Body_y[628] = c_Body_y[627];
                    end else begin
                        n_Body_x[628] = c_Body_x[c_Size-1];
                        n_Body_y[628] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 629) begin
                        n_Body_x[629] = c_Body_x[628];
                        n_Body_y[629] = c_Body_y[628];
                    end else begin
                        n_Body_x[629] = c_Body_x[c_Size-1];
                        n_Body_y[629] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 630) begin
                        n_Body_x[630] = c_Body_x[629];
                        n_Body_y[630] = c_Body_y[629];
                    end else begin
                        n_Body_x[630] = c_Body_x[c_Size-1];
                        n_Body_y[630] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 631) begin
                        n_Body_x[631] = c_Body_x[630];
                        n_Body_y[631] = c_Body_y[630];
                    end else begin
                        n_Body_x[631] = c_Body_x[c_Size-1];
                        n_Body_y[631] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 632) begin
                        n_Body_x[632] = c_Body_x[631];
                        n_Body_y[632] = c_Body_y[631];
                    end else begin
                        n_Body_x[632] = c_Body_x[c_Size-1];
                        n_Body_y[632] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 633) begin
                        n_Body_x[633] = c_Body_x[632];
                        n_Body_y[633] = c_Body_y[632];
                    end else begin
                        n_Body_x[633] = c_Body_x[c_Size-1];
                        n_Body_y[633] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 634) begin
                        n_Body_x[634] = c_Body_x[633];
                        n_Body_y[634] = c_Body_y[633];
                    end else begin
                        n_Body_x[634] = c_Body_x[c_Size-1];
                        n_Body_y[634] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 635) begin
                        n_Body_x[635] = c_Body_x[634];
                        n_Body_y[635] = c_Body_y[634];
                    end else begin
                        n_Body_x[635] = c_Body_x[c_Size-1];
                        n_Body_y[635] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 636) begin
                        n_Body_x[636] = c_Body_x[635];
                        n_Body_y[636] = c_Body_y[635];
                    end else begin
                        n_Body_x[636] = c_Body_x[c_Size-1];
                        n_Body_y[636] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 637) begin
                        n_Body_x[637] = c_Body_x[636];
                        n_Body_y[637] = c_Body_y[636];
                    end else begin
                        n_Body_x[637] = c_Body_x[c_Size-1];
                        n_Body_y[637] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 638) begin
                        n_Body_x[638] = c_Body_x[637];
                        n_Body_y[638] = c_Body_y[637];
                    end else begin
                        n_Body_x[638] = c_Body_x[c_Size-1];
                        n_Body_y[638] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 639) begin
                        n_Body_x[639] = c_Body_x[638];
                        n_Body_y[639] = c_Body_y[638];
                    end else begin
                        n_Body_x[639] = c_Body_x[c_Size-1];
                        n_Body_y[639] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 640) begin
                        n_Body_x[640] = c_Body_x[639];
                        n_Body_y[640] = c_Body_y[639];
                    end else begin
                        n_Body_x[640] = c_Body_x[c_Size-1];
                        n_Body_y[640] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 641) begin
                        n_Body_x[641] = c_Body_x[640];
                        n_Body_y[641] = c_Body_y[640];
                    end else begin
                        n_Body_x[641] = c_Body_x[c_Size-1];
                        n_Body_y[641] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 642) begin
                        n_Body_x[642] = c_Body_x[641];
                        n_Body_y[642] = c_Body_y[641];
                    end else begin
                        n_Body_x[642] = c_Body_x[c_Size-1];
                        n_Body_y[642] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 643) begin
                        n_Body_x[643] = c_Body_x[642];
                        n_Body_y[643] = c_Body_y[642];
                    end else begin
                        n_Body_x[643] = c_Body_x[c_Size-1];
                        n_Body_y[643] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 644) begin
                        n_Body_x[644] = c_Body_x[643];
                        n_Body_y[644] = c_Body_y[643];
                    end else begin
                        n_Body_x[644] = c_Body_x[c_Size-1];
                        n_Body_y[644] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 645) begin
                        n_Body_x[645] = c_Body_x[644];
                        n_Body_y[645] = c_Body_y[644];
                    end else begin
                        n_Body_x[645] = c_Body_x[c_Size-1];
                        n_Body_y[645] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 646) begin
                        n_Body_x[646] = c_Body_x[645];
                        n_Body_y[646] = c_Body_y[645];
                    end else begin
                        n_Body_x[646] = c_Body_x[c_Size-1];
                        n_Body_y[646] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 647) begin
                        n_Body_x[647] = c_Body_x[646];
                        n_Body_y[647] = c_Body_y[646];
                    end else begin
                        n_Body_x[647] = c_Body_x[c_Size-1];
                        n_Body_y[647] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 648) begin
                        n_Body_x[648] = c_Body_x[647];
                        n_Body_y[648] = c_Body_y[647];
                    end else begin
                        n_Body_x[648] = c_Body_x[c_Size-1];
                        n_Body_y[648] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 649) begin
                        n_Body_x[649] = c_Body_x[648];
                        n_Body_y[649] = c_Body_y[648];
                    end else begin
                        n_Body_x[649] = c_Body_x[c_Size-1];
                        n_Body_y[649] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 650) begin
                        n_Body_x[650] = c_Body_x[649];
                        n_Body_y[650] = c_Body_y[649];
                    end else begin
                        n_Body_x[650] = c_Body_x[c_Size-1];
                        n_Body_y[650] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 651) begin
                        n_Body_x[651] = c_Body_x[650];
                        n_Body_y[651] = c_Body_y[650];
                    end else begin
                        n_Body_x[651] = c_Body_x[c_Size-1];
                        n_Body_y[651] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 652) begin
                        n_Body_x[652] = c_Body_x[651];
                        n_Body_y[652] = c_Body_y[651];
                    end else begin
                        n_Body_x[652] = c_Body_x[c_Size-1];
                        n_Body_y[652] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 653) begin
                        n_Body_x[653] = c_Body_x[652];
                        n_Body_y[653] = c_Body_y[652];
                    end else begin
                        n_Body_x[653] = c_Body_x[c_Size-1];
                        n_Body_y[653] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 654) begin
                        n_Body_x[654] = c_Body_x[653];
                        n_Body_y[654] = c_Body_y[653];
                    end else begin
                        n_Body_x[654] = c_Body_x[c_Size-1];
                        n_Body_y[654] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 655) begin
                        n_Body_x[655] = c_Body_x[654];
                        n_Body_y[655] = c_Body_y[654];
                    end else begin
                        n_Body_x[655] = c_Body_x[c_Size-1];
                        n_Body_y[655] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 656) begin
                        n_Body_x[656] = c_Body_x[655];
                        n_Body_y[656] = c_Body_y[655];
                    end else begin
                        n_Body_x[656] = c_Body_x[c_Size-1];
                        n_Body_y[656] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 657) begin
                        n_Body_x[657] = c_Body_x[656];
                        n_Body_y[657] = c_Body_y[656];
                    end else begin
                        n_Body_x[657] = c_Body_x[c_Size-1];
                        n_Body_y[657] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 658) begin
                        n_Body_x[658] = c_Body_x[657];
                        n_Body_y[658] = c_Body_y[657];
                    end else begin
                        n_Body_x[658] = c_Body_x[c_Size-1];
                        n_Body_y[658] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 659) begin
                        n_Body_x[659] = c_Body_x[658];
                        n_Body_y[659] = c_Body_y[658];
                    end else begin
                        n_Body_x[659] = c_Body_x[c_Size-1];
                        n_Body_y[659] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 660) begin
                        n_Body_x[660] = c_Body_x[659];
                        n_Body_y[660] = c_Body_y[659];
                    end else begin
                        n_Body_x[660] = c_Body_x[c_Size-1];
                        n_Body_y[660] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 661) begin
                        n_Body_x[661] = c_Body_x[660];
                        n_Body_y[661] = c_Body_y[660];
                    end else begin
                        n_Body_x[661] = c_Body_x[c_Size-1];
                        n_Body_y[661] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 662) begin
                        n_Body_x[662] = c_Body_x[661];
                        n_Body_y[662] = c_Body_y[661];
                    end else begin
                        n_Body_x[662] = c_Body_x[c_Size-1];
                        n_Body_y[662] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 663) begin
                        n_Body_x[663] = c_Body_x[662];
                        n_Body_y[663] = c_Body_y[662];
                    end else begin
                        n_Body_x[663] = c_Body_x[c_Size-1];
                        n_Body_y[663] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 664) begin
                        n_Body_x[664] = c_Body_x[663];
                        n_Body_y[664] = c_Body_y[663];
                    end else begin
                        n_Body_x[664] = c_Body_x[c_Size-1];
                        n_Body_y[664] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 665) begin
                        n_Body_x[665] = c_Body_x[664];
                        n_Body_y[665] = c_Body_y[664];
                    end else begin
                        n_Body_x[665] = c_Body_x[c_Size-1];
                        n_Body_y[665] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 666) begin
                        n_Body_x[666] = c_Body_x[665];
                        n_Body_y[666] = c_Body_y[665];
                    end else begin
                        n_Body_x[666] = c_Body_x[c_Size-1];
                        n_Body_y[666] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 667) begin
                        n_Body_x[667] = c_Body_x[666];
                        n_Body_y[667] = c_Body_y[666];
                    end else begin
                        n_Body_x[667] = c_Body_x[c_Size-1];
                        n_Body_y[667] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 668) begin
                        n_Body_x[668] = c_Body_x[667];
                        n_Body_y[668] = c_Body_y[667];
                    end else begin
                        n_Body_x[668] = c_Body_x[c_Size-1];
                        n_Body_y[668] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 669) begin
                        n_Body_x[669] = c_Body_x[668];
                        n_Body_y[669] = c_Body_y[668];
                    end else begin
                        n_Body_x[669] = c_Body_x[c_Size-1];
                        n_Body_y[669] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 670) begin
                        n_Body_x[670] = c_Body_x[669];
                        n_Body_y[670] = c_Body_y[669];
                    end else begin
                        n_Body_x[670] = c_Body_x[c_Size-1];
                        n_Body_y[670] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 671) begin
                        n_Body_x[671] = c_Body_x[670];
                        n_Body_y[671] = c_Body_y[670];
                    end else begin
                        n_Body_x[671] = c_Body_x[c_Size-1];
                        n_Body_y[671] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 672) begin
                        n_Body_x[672] = c_Body_x[671];
                        n_Body_y[672] = c_Body_y[671];
                    end else begin
                        n_Body_x[672] = c_Body_x[c_Size-1];
                        n_Body_y[672] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 673) begin
                        n_Body_x[673] = c_Body_x[672];
                        n_Body_y[673] = c_Body_y[672];
                    end else begin
                        n_Body_x[673] = c_Body_x[c_Size-1];
                        n_Body_y[673] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 674) begin
                        n_Body_x[674] = c_Body_x[673];
                        n_Body_y[674] = c_Body_y[673];
                    end else begin
                        n_Body_x[674] = c_Body_x[c_Size-1];
                        n_Body_y[674] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 675) begin
                        n_Body_x[675] = c_Body_x[674];
                        n_Body_y[675] = c_Body_y[674];
                    end else begin
                        n_Body_x[675] = c_Body_x[c_Size-1];
                        n_Body_y[675] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 676) begin
                        n_Body_x[676] = c_Body_x[675];
                        n_Body_y[676] = c_Body_y[675];
                    end else begin
                        n_Body_x[676] = c_Body_x[c_Size-1];
                        n_Body_y[676] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 677) begin
                        n_Body_x[677] = c_Body_x[676];
                        n_Body_y[677] = c_Body_y[676];
                    end else begin
                        n_Body_x[677] = c_Body_x[c_Size-1];
                        n_Body_y[677] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 678) begin
                        n_Body_x[678] = c_Body_x[677];
                        n_Body_y[678] = c_Body_y[677];
                    end else begin
                        n_Body_x[678] = c_Body_x[c_Size-1];
                        n_Body_y[678] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 679) begin
                        n_Body_x[679] = c_Body_x[678];
                        n_Body_y[679] = c_Body_y[678];
                    end else begin
                        n_Body_x[679] = c_Body_x[c_Size-1];
                        n_Body_y[679] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 680) begin
                        n_Body_x[680] = c_Body_x[679];
                        n_Body_y[680] = c_Body_y[679];
                    end else begin
                        n_Body_x[680] = c_Body_x[c_Size-1];
                        n_Body_y[680] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 681) begin
                        n_Body_x[681] = c_Body_x[680];
                        n_Body_y[681] = c_Body_y[680];
                    end else begin
                        n_Body_x[681] = c_Body_x[c_Size-1];
                        n_Body_y[681] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 682) begin
                        n_Body_x[682] = c_Body_x[681];
                        n_Body_y[682] = c_Body_y[681];
                    end else begin
                        n_Body_x[682] = c_Body_x[c_Size-1];
                        n_Body_y[682] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 683) begin
                        n_Body_x[683] = c_Body_x[682];
                        n_Body_y[683] = c_Body_y[682];
                    end else begin
                        n_Body_x[683] = c_Body_x[c_Size-1];
                        n_Body_y[683] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 684) begin
                        n_Body_x[684] = c_Body_x[683];
                        n_Body_y[684] = c_Body_y[683];
                    end else begin
                        n_Body_x[684] = c_Body_x[c_Size-1];
                        n_Body_y[684] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 685) begin
                        n_Body_x[685] = c_Body_x[684];
                        n_Body_y[685] = c_Body_y[684];
                    end else begin
                        n_Body_x[685] = c_Body_x[c_Size-1];
                        n_Body_y[685] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 686) begin
                        n_Body_x[686] = c_Body_x[685];
                        n_Body_y[686] = c_Body_y[685];
                    end else begin
                        n_Body_x[686] = c_Body_x[c_Size-1];
                        n_Body_y[686] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 687) begin
                        n_Body_x[687] = c_Body_x[686];
                        n_Body_y[687] = c_Body_y[686];
                    end else begin
                        n_Body_x[687] = c_Body_x[c_Size-1];
                        n_Body_y[687] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 688) begin
                        n_Body_x[688] = c_Body_x[687];
                        n_Body_y[688] = c_Body_y[687];
                    end else begin
                        n_Body_x[688] = c_Body_x[c_Size-1];
                        n_Body_y[688] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 689) begin
                        n_Body_x[689] = c_Body_x[688];
                        n_Body_y[689] = c_Body_y[688];
                    end else begin
                        n_Body_x[689] = c_Body_x[c_Size-1];
                        n_Body_y[689] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 690) begin
                        n_Body_x[690] = c_Body_x[689];
                        n_Body_y[690] = c_Body_y[689];
                    end else begin
                        n_Body_x[690] = c_Body_x[c_Size-1];
                        n_Body_y[690] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 691) begin
                        n_Body_x[691] = c_Body_x[690];
                        n_Body_y[691] = c_Body_y[690];
                    end else begin
                        n_Body_x[691] = c_Body_x[c_Size-1];
                        n_Body_y[691] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 692) begin
                        n_Body_x[692] = c_Body_x[691];
                        n_Body_y[692] = c_Body_y[691];
                    end else begin
                        n_Body_x[692] = c_Body_x[c_Size-1];
                        n_Body_y[692] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 693) begin
                        n_Body_x[693] = c_Body_x[692];
                        n_Body_y[693] = c_Body_y[692];
                    end else begin
                        n_Body_x[693] = c_Body_x[c_Size-1];
                        n_Body_y[693] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 694) begin
                        n_Body_x[694] = c_Body_x[693];
                        n_Body_y[694] = c_Body_y[693];
                    end else begin
                        n_Body_x[694] = c_Body_x[c_Size-1];
                        n_Body_y[694] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 695) begin
                        n_Body_x[695] = c_Body_x[694];
                        n_Body_y[695] = c_Body_y[694];
                    end else begin
                        n_Body_x[695] = c_Body_x[c_Size-1];
                        n_Body_y[695] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 696) begin
                        n_Body_x[696] = c_Body_x[695];
                        n_Body_y[696] = c_Body_y[695];
                    end else begin
                        n_Body_x[696] = c_Body_x[c_Size-1];
                        n_Body_y[696] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 697) begin
                        n_Body_x[697] = c_Body_x[696];
                        n_Body_y[697] = c_Body_y[696];
                    end else begin
                        n_Body_x[697] = c_Body_x[c_Size-1];
                        n_Body_y[697] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 698) begin
                        n_Body_x[698] = c_Body_x[697];
                        n_Body_y[698] = c_Body_y[697];
                    end else begin
                        n_Body_x[698] = c_Body_x[c_Size-1];
                        n_Body_y[698] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 699) begin
                        n_Body_x[699] = c_Body_x[698];
                        n_Body_y[699] = c_Body_y[698];
                    end else begin
                        n_Body_x[699] = c_Body_x[c_Size-1];
                        n_Body_y[699] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 700) begin
                        n_Body_x[700] = c_Body_x[699];
                        n_Body_y[700] = c_Body_y[699];
                    end else begin
                        n_Body_x[700] = c_Body_x[c_Size-1];
                        n_Body_y[700] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 701) begin
                        n_Body_x[701] = c_Body_x[700];
                        n_Body_y[701] = c_Body_y[700];
                    end else begin
                        n_Body_x[701] = c_Body_x[c_Size-1];
                        n_Body_y[701] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 702) begin
                        n_Body_x[702] = c_Body_x[701];
                        n_Body_y[702] = c_Body_y[701];
                    end else begin
                        n_Body_x[702] = c_Body_x[c_Size-1];
                        n_Body_y[702] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 703) begin
                        n_Body_x[703] = c_Body_x[702];
                        n_Body_y[703] = c_Body_y[702];
                    end else begin
                        n_Body_x[703] = c_Body_x[c_Size-1];
                        n_Body_y[703] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 704) begin
                        n_Body_x[704] = c_Body_x[703];
                        n_Body_y[704] = c_Body_y[703];
                    end else begin
                        n_Body_x[704] = c_Body_x[c_Size-1];
                        n_Body_y[704] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 705) begin
                        n_Body_x[705] = c_Body_x[704];
                        n_Body_y[705] = c_Body_y[704];
                    end else begin
                        n_Body_x[705] = c_Body_x[c_Size-1];
                        n_Body_y[705] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 706) begin
                        n_Body_x[706] = c_Body_x[705];
                        n_Body_y[706] = c_Body_y[705];
                    end else begin
                        n_Body_x[706] = c_Body_x[c_Size-1];
                        n_Body_y[706] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 707) begin
                        n_Body_x[707] = c_Body_x[706];
                        n_Body_y[707] = c_Body_y[706];
                    end else begin
                        n_Body_x[707] = c_Body_x[c_Size-1];
                        n_Body_y[707] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 708) begin
                        n_Body_x[708] = c_Body_x[707];
                        n_Body_y[708] = c_Body_y[707];
                    end else begin
                        n_Body_x[708] = c_Body_x[c_Size-1];
                        n_Body_y[708] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 709) begin
                        n_Body_x[709] = c_Body_x[708];
                        n_Body_y[709] = c_Body_y[708];
                    end else begin
                        n_Body_x[709] = c_Body_x[c_Size-1];
                        n_Body_y[709] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 710) begin
                        n_Body_x[710] = c_Body_x[709];
                        n_Body_y[710] = c_Body_y[709];
                    end else begin
                        n_Body_x[710] = c_Body_x[c_Size-1];
                        n_Body_y[710] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 711) begin
                        n_Body_x[711] = c_Body_x[710];
                        n_Body_y[711] = c_Body_y[710];
                    end else begin
                        n_Body_x[711] = c_Body_x[c_Size-1];
                        n_Body_y[711] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 712) begin
                        n_Body_x[712] = c_Body_x[711];
                        n_Body_y[712] = c_Body_y[711];
                    end else begin
                        n_Body_x[712] = c_Body_x[c_Size-1];
                        n_Body_y[712] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 713) begin
                        n_Body_x[713] = c_Body_x[712];
                        n_Body_y[713] = c_Body_y[712];
                    end else begin
                        n_Body_x[713] = c_Body_x[c_Size-1];
                        n_Body_y[713] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 714) begin
                        n_Body_x[714] = c_Body_x[713];
                        n_Body_y[714] = c_Body_y[713];
                    end else begin
                        n_Body_x[714] = c_Body_x[c_Size-1];
                        n_Body_y[714] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 715) begin
                        n_Body_x[715] = c_Body_x[714];
                        n_Body_y[715] = c_Body_y[714];
                    end else begin
                        n_Body_x[715] = c_Body_x[c_Size-1];
                        n_Body_y[715] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 716) begin
                        n_Body_x[716] = c_Body_x[715];
                        n_Body_y[716] = c_Body_y[715];
                    end else begin
                        n_Body_x[716] = c_Body_x[c_Size-1];
                        n_Body_y[716] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 717) begin
                        n_Body_x[717] = c_Body_x[716];
                        n_Body_y[717] = c_Body_y[716];
                    end else begin
                        n_Body_x[717] = c_Body_x[c_Size-1];
                        n_Body_y[717] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 718) begin
                        n_Body_x[718] = c_Body_x[717];
                        n_Body_y[718] = c_Body_y[717];
                    end else begin
                        n_Body_x[718] = c_Body_x[c_Size-1];
                        n_Body_y[718] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 719) begin
                        n_Body_x[719] = c_Body_x[718];
                        n_Body_y[719] = c_Body_y[718];
                    end else begin
                        n_Body_x[719] = c_Body_x[c_Size-1];
                        n_Body_y[719] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 720) begin
                        n_Body_x[720] = c_Body_x[719];
                        n_Body_y[720] = c_Body_y[719];
                    end else begin
                        n_Body_x[720] = c_Body_x[c_Size-1];
                        n_Body_y[720] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 721) begin
                        n_Body_x[721] = c_Body_x[720];
                        n_Body_y[721] = c_Body_y[720];
                    end else begin
                        n_Body_x[721] = c_Body_x[c_Size-1];
                        n_Body_y[721] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 722) begin
                        n_Body_x[722] = c_Body_x[721];
                        n_Body_y[722] = c_Body_y[721];
                    end else begin
                        n_Body_x[722] = c_Body_x[c_Size-1];
                        n_Body_y[722] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 723) begin
                        n_Body_x[723] = c_Body_x[722];
                        n_Body_y[723] = c_Body_y[722];
                    end else begin
                        n_Body_x[723] = c_Body_x[c_Size-1];
                        n_Body_y[723] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 724) begin
                        n_Body_x[724] = c_Body_x[723];
                        n_Body_y[724] = c_Body_y[723];
                    end else begin
                        n_Body_x[724] = c_Body_x[c_Size-1];
                        n_Body_y[724] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 725) begin
                        n_Body_x[725] = c_Body_x[724];
                        n_Body_y[725] = c_Body_y[724];
                    end else begin
                        n_Body_x[725] = c_Body_x[c_Size-1];
                        n_Body_y[725] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 726) begin
                        n_Body_x[726] = c_Body_x[725];
                        n_Body_y[726] = c_Body_y[725];
                    end else begin
                        n_Body_x[726] = c_Body_x[c_Size-1];
                        n_Body_y[726] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 727) begin
                        n_Body_x[727] = c_Body_x[726];
                        n_Body_y[727] = c_Body_y[726];
                    end else begin
                        n_Body_x[727] = c_Body_x[c_Size-1];
                        n_Body_y[727] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 728) begin
                        n_Body_x[728] = c_Body_x[727];
                        n_Body_y[728] = c_Body_y[727];
                    end else begin
                        n_Body_x[728] = c_Body_x[c_Size-1];
                        n_Body_y[728] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 729) begin
                        n_Body_x[729] = c_Body_x[728];
                        n_Body_y[729] = c_Body_y[728];
                    end else begin
                        n_Body_x[729] = c_Body_x[c_Size-1];
                        n_Body_y[729] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 730) begin
                        n_Body_x[730] = c_Body_x[729];
                        n_Body_y[730] = c_Body_y[729];
                    end else begin
                        n_Body_x[730] = c_Body_x[c_Size-1];
                        n_Body_y[730] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 731) begin
                        n_Body_x[731] = c_Body_x[730];
                        n_Body_y[731] = c_Body_y[730];
                    end else begin
                        n_Body_x[731] = c_Body_x[c_Size-1];
                        n_Body_y[731] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 732) begin
                        n_Body_x[732] = c_Body_x[731];
                        n_Body_y[732] = c_Body_y[731];
                    end else begin
                        n_Body_x[732] = c_Body_x[c_Size-1];
                        n_Body_y[732] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 733) begin
                        n_Body_x[733] = c_Body_x[732];
                        n_Body_y[733] = c_Body_y[732];
                    end else begin
                        n_Body_x[733] = c_Body_x[c_Size-1];
                        n_Body_y[733] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 734) begin
                        n_Body_x[734] = c_Body_x[733];
                        n_Body_y[734] = c_Body_y[733];
                    end else begin
                        n_Body_x[734] = c_Body_x[c_Size-1];
                        n_Body_y[734] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 735) begin
                        n_Body_x[735] = c_Body_x[734];
                        n_Body_y[735] = c_Body_y[734];
                    end else begin
                        n_Body_x[735] = c_Body_x[c_Size-1];
                        n_Body_y[735] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 736) begin
                        n_Body_x[736] = c_Body_x[735];
                        n_Body_y[736] = c_Body_y[735];
                    end else begin
                        n_Body_x[736] = c_Body_x[c_Size-1];
                        n_Body_y[736] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 737) begin
                        n_Body_x[737] = c_Body_x[736];
                        n_Body_y[737] = c_Body_y[736];
                    end else begin
                        n_Body_x[737] = c_Body_x[c_Size-1];
                        n_Body_y[737] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 738) begin
                        n_Body_x[738] = c_Body_x[737];
                        n_Body_y[738] = c_Body_y[737];
                    end else begin
                        n_Body_x[738] = c_Body_x[c_Size-1];
                        n_Body_y[738] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 739) begin
                        n_Body_x[739] = c_Body_x[738];
                        n_Body_y[739] = c_Body_y[738];
                    end else begin
                        n_Body_x[739] = c_Body_x[c_Size-1];
                        n_Body_y[739] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 740) begin
                        n_Body_x[740] = c_Body_x[739];
                        n_Body_y[740] = c_Body_y[739];
                    end else begin
                        n_Body_x[740] = c_Body_x[c_Size-1];
                        n_Body_y[740] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 741) begin
                        n_Body_x[741] = c_Body_x[740];
                        n_Body_y[741] = c_Body_y[740];
                    end else begin
                        n_Body_x[741] = c_Body_x[c_Size-1];
                        n_Body_y[741] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 742) begin
                        n_Body_x[742] = c_Body_x[741];
                        n_Body_y[742] = c_Body_y[741];
                    end else begin
                        n_Body_x[742] = c_Body_x[c_Size-1];
                        n_Body_y[742] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 743) begin
                        n_Body_x[743] = c_Body_x[742];
                        n_Body_y[743] = c_Body_y[742];
                    end else begin
                        n_Body_x[743] = c_Body_x[c_Size-1];
                        n_Body_y[743] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 744) begin
                        n_Body_x[744] = c_Body_x[743];
                        n_Body_y[744] = c_Body_y[743];
                    end else begin
                        n_Body_x[744] = c_Body_x[c_Size-1];
                        n_Body_y[744] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 745) begin
                        n_Body_x[745] = c_Body_x[744];
                        n_Body_y[745] = c_Body_y[744];
                    end else begin
                        n_Body_x[745] = c_Body_x[c_Size-1];
                        n_Body_y[745] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 746) begin
                        n_Body_x[746] = c_Body_x[745];
                        n_Body_y[746] = c_Body_y[745];
                    end else begin
                        n_Body_x[746] = c_Body_x[c_Size-1];
                        n_Body_y[746] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 747) begin
                        n_Body_x[747] = c_Body_x[746];
                        n_Body_y[747] = c_Body_y[746];
                    end else begin
                        n_Body_x[747] = c_Body_x[c_Size-1];
                        n_Body_y[747] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 748) begin
                        n_Body_x[748] = c_Body_x[747];
                        n_Body_y[748] = c_Body_y[747];
                    end else begin
                        n_Body_x[748] = c_Body_x[c_Size-1];
                        n_Body_y[748] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 749) begin
                        n_Body_x[749] = c_Body_x[748];
                        n_Body_y[749] = c_Body_y[748];
                    end else begin
                        n_Body_x[749] = c_Body_x[c_Size-1];
                        n_Body_y[749] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 750) begin
                        n_Body_x[750] = c_Body_x[749];
                        n_Body_y[750] = c_Body_y[749];
                    end else begin
                        n_Body_x[750] = c_Body_x[c_Size-1];
                        n_Body_y[750] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 751) begin
                        n_Body_x[751] = c_Body_x[750];
                        n_Body_y[751] = c_Body_y[750];
                    end else begin
                        n_Body_x[751] = c_Body_x[c_Size-1];
                        n_Body_y[751] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 752) begin
                        n_Body_x[752] = c_Body_x[751];
                        n_Body_y[752] = c_Body_y[751];
                    end else begin
                        n_Body_x[752] = c_Body_x[c_Size-1];
                        n_Body_y[752] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 753) begin
                        n_Body_x[753] = c_Body_x[752];
                        n_Body_y[753] = c_Body_y[752];
                    end else begin
                        n_Body_x[753] = c_Body_x[c_Size-1];
                        n_Body_y[753] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 754) begin
                        n_Body_x[754] = c_Body_x[753];
                        n_Body_y[754] = c_Body_y[753];
                    end else begin
                        n_Body_x[754] = c_Body_x[c_Size-1];
                        n_Body_y[754] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 755) begin
                        n_Body_x[755] = c_Body_x[754];
                        n_Body_y[755] = c_Body_y[754];
                    end else begin
                        n_Body_x[755] = c_Body_x[c_Size-1];
                        n_Body_y[755] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 756) begin
                        n_Body_x[756] = c_Body_x[755];
                        n_Body_y[756] = c_Body_y[755];
                    end else begin
                        n_Body_x[756] = c_Body_x[c_Size-1];
                        n_Body_y[756] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 757) begin
                        n_Body_x[757] = c_Body_x[756];
                        n_Body_y[757] = c_Body_y[756];
                    end else begin
                        n_Body_x[757] = c_Body_x[c_Size-1];
                        n_Body_y[757] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 758) begin
                        n_Body_x[758] = c_Body_x[757];
                        n_Body_y[758] = c_Body_y[757];
                    end else begin
                        n_Body_x[758] = c_Body_x[c_Size-1];
                        n_Body_y[758] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 759) begin
                        n_Body_x[759] = c_Body_x[758];
                        n_Body_y[759] = c_Body_y[758];
                    end else begin
                        n_Body_x[759] = c_Body_x[c_Size-1];
                        n_Body_y[759] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 760) begin
                        n_Body_x[760] = c_Body_x[759];
                        n_Body_y[760] = c_Body_y[759];
                    end else begin
                        n_Body_x[760] = c_Body_x[c_Size-1];
                        n_Body_y[760] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 761) begin
                        n_Body_x[761] = c_Body_x[760];
                        n_Body_y[761] = c_Body_y[760];
                    end else begin
                        n_Body_x[761] = c_Body_x[c_Size-1];
                        n_Body_y[761] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 762) begin
                        n_Body_x[762] = c_Body_x[761];
                        n_Body_y[762] = c_Body_y[761];
                    end else begin
                        n_Body_x[762] = c_Body_x[c_Size-1];
                        n_Body_y[762] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 763) begin
                        n_Body_x[763] = c_Body_x[762];
                        n_Body_y[763] = c_Body_y[762];
                    end else begin
                        n_Body_x[763] = c_Body_x[c_Size-1];
                        n_Body_y[763] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 764) begin
                        n_Body_x[764] = c_Body_x[763];
                        n_Body_y[764] = c_Body_y[763];
                    end else begin
                        n_Body_x[764] = c_Body_x[c_Size-1];
                        n_Body_y[764] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 765) begin
                        n_Body_x[765] = c_Body_x[764];
                        n_Body_y[765] = c_Body_y[764];
                    end else begin
                        n_Body_x[765] = c_Body_x[c_Size-1];
                        n_Body_y[765] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 766) begin
                        n_Body_x[766] = c_Body_x[765];
                        n_Body_y[766] = c_Body_y[765];
                    end else begin
                        n_Body_x[766] = c_Body_x[c_Size-1];
                        n_Body_y[766] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 767) begin
                        n_Body_x[767] = c_Body_x[766];
                        n_Body_y[767] = c_Body_y[766];
                    end else begin
                        n_Body_x[767] = c_Body_x[c_Size-1];
                        n_Body_y[767] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 768) begin
                        n_Body_x[768] = c_Body_x[767];
                        n_Body_y[768] = c_Body_y[767];
                    end else begin
                        n_Body_x[768] = c_Body_x[c_Size-1];
                        n_Body_y[768] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 769) begin
                        n_Body_x[769] = c_Body_x[768];
                        n_Body_y[769] = c_Body_y[768];
                    end else begin
                        n_Body_x[769] = c_Body_x[c_Size-1];
                        n_Body_y[769] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 770) begin
                        n_Body_x[770] = c_Body_x[769];
                        n_Body_y[770] = c_Body_y[769];
                    end else begin
                        n_Body_x[770] = c_Body_x[c_Size-1];
                        n_Body_y[770] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 771) begin
                        n_Body_x[771] = c_Body_x[770];
                        n_Body_y[771] = c_Body_y[770];
                    end else begin
                        n_Body_x[771] = c_Body_x[c_Size-1];
                        n_Body_y[771] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 772) begin
                        n_Body_x[772] = c_Body_x[771];
                        n_Body_y[772] = c_Body_y[771];
                    end else begin
                        n_Body_x[772] = c_Body_x[c_Size-1];
                        n_Body_y[772] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 773) begin
                        n_Body_x[773] = c_Body_x[772];
                        n_Body_y[773] = c_Body_y[772];
                    end else begin
                        n_Body_x[773] = c_Body_x[c_Size-1];
                        n_Body_y[773] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 774) begin
                        n_Body_x[774] = c_Body_x[773];
                        n_Body_y[774] = c_Body_y[773];
                    end else begin
                        n_Body_x[774] = c_Body_x[c_Size-1];
                        n_Body_y[774] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 775) begin
                        n_Body_x[775] = c_Body_x[774];
                        n_Body_y[775] = c_Body_y[774];
                    end else begin
                        n_Body_x[775] = c_Body_x[c_Size-1];
                        n_Body_y[775] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 776) begin
                        n_Body_x[776] = c_Body_x[775];
                        n_Body_y[776] = c_Body_y[775];
                    end else begin
                        n_Body_x[776] = c_Body_x[c_Size-1];
                        n_Body_y[776] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 777) begin
                        n_Body_x[777] = c_Body_x[776];
                        n_Body_y[777] = c_Body_y[776];
                    end else begin
                        n_Body_x[777] = c_Body_x[c_Size-1];
                        n_Body_y[777] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 778) begin
                        n_Body_x[778] = c_Body_x[777];
                        n_Body_y[778] = c_Body_y[777];
                    end else begin
                        n_Body_x[778] = c_Body_x[c_Size-1];
                        n_Body_y[778] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 779) begin
                        n_Body_x[779] = c_Body_x[778];
                        n_Body_y[779] = c_Body_y[778];
                    end else begin
                        n_Body_x[779] = c_Body_x[c_Size-1];
                        n_Body_y[779] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 780) begin
                        n_Body_x[780] = c_Body_x[779];
                        n_Body_y[780] = c_Body_y[779];
                    end else begin
                        n_Body_x[780] = c_Body_x[c_Size-1];
                        n_Body_y[780] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 781) begin
                        n_Body_x[781] = c_Body_x[780];
                        n_Body_y[781] = c_Body_y[780];
                    end else begin
                        n_Body_x[781] = c_Body_x[c_Size-1];
                        n_Body_y[781] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 782) begin
                        n_Body_x[782] = c_Body_x[781];
                        n_Body_y[782] = c_Body_y[781];
                    end else begin
                        n_Body_x[782] = c_Body_x[c_Size-1];
                        n_Body_y[782] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 783) begin
                        n_Body_x[783] = c_Body_x[782];
                        n_Body_y[783] = c_Body_y[782];
                    end else begin
                        n_Body_x[783] = c_Body_x[c_Size-1];
                        n_Body_y[783] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 784) begin
                        n_Body_x[784] = c_Body_x[783];
                        n_Body_y[784] = c_Body_y[783];
                    end else begin
                        n_Body_x[784] = c_Body_x[c_Size-1];
                        n_Body_y[784] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 785) begin
                        n_Body_x[785] = c_Body_x[784];
                        n_Body_y[785] = c_Body_y[784];
                    end else begin
                        n_Body_x[785] = c_Body_x[c_Size-1];
                        n_Body_y[785] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 786) begin
                        n_Body_x[786] = c_Body_x[785];
                        n_Body_y[786] = c_Body_y[785];
                    end else begin
                        n_Body_x[786] = c_Body_x[c_Size-1];
                        n_Body_y[786] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 787) begin
                        n_Body_x[787] = c_Body_x[786];
                        n_Body_y[787] = c_Body_y[786];
                    end else begin
                        n_Body_x[787] = c_Body_x[c_Size-1];
                        n_Body_y[787] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 788) begin
                        n_Body_x[788] = c_Body_x[787];
                        n_Body_y[788] = c_Body_y[787];
                    end else begin
                        n_Body_x[788] = c_Body_x[c_Size-1];
                        n_Body_y[788] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 789) begin
                        n_Body_x[789] = c_Body_x[788];
                        n_Body_y[789] = c_Body_y[788];
                    end else begin
                        n_Body_x[789] = c_Body_x[c_Size-1];
                        n_Body_y[789] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 790) begin
                        n_Body_x[790] = c_Body_x[789];
                        n_Body_y[790] = c_Body_y[789];
                    end else begin
                        n_Body_x[790] = c_Body_x[c_Size-1];
                        n_Body_y[790] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 791) begin
                        n_Body_x[791] = c_Body_x[790];
                        n_Body_y[791] = c_Body_y[790];
                    end else begin
                        n_Body_x[791] = c_Body_x[c_Size-1];
                        n_Body_y[791] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 792) begin
                        n_Body_x[792] = c_Body_x[791];
                        n_Body_y[792] = c_Body_y[791];
                    end else begin
                        n_Body_x[792] = c_Body_x[c_Size-1];
                        n_Body_y[792] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 793) begin
                        n_Body_x[793] = c_Body_x[792];
                        n_Body_y[793] = c_Body_y[792];
                    end else begin
                        n_Body_x[793] = c_Body_x[c_Size-1];
                        n_Body_y[793] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 794) begin
                        n_Body_x[794] = c_Body_x[793];
                        n_Body_y[794] = c_Body_y[793];
                    end else begin
                        n_Body_x[794] = c_Body_x[c_Size-1];
                        n_Body_y[794] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 795) begin
                        n_Body_x[795] = c_Body_x[794];
                        n_Body_y[795] = c_Body_y[794];
                    end else begin
                        n_Body_x[795] = c_Body_x[c_Size-1];
                        n_Body_y[795] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 796) begin
                        n_Body_x[796] = c_Body_x[795];
                        n_Body_y[796] = c_Body_y[795];
                    end else begin
                        n_Body_x[796] = c_Body_x[c_Size-1];
                        n_Body_y[796] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 797) begin
                        n_Body_x[797] = c_Body_x[796];
                        n_Body_y[797] = c_Body_y[796];
                    end else begin
                        n_Body_x[797] = c_Body_x[c_Size-1];
                        n_Body_y[797] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 798) begin
                        n_Body_x[798] = c_Body_x[797];
                        n_Body_y[798] = c_Body_y[797];
                    end else begin
                        n_Body_x[798] = c_Body_x[c_Size-1];
                        n_Body_y[798] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 799) begin
                        n_Body_x[799] = c_Body_x[798];
                        n_Body_y[799] = c_Body_y[798];
                    end else begin
                        n_Body_x[799] = c_Body_x[c_Size-1];
                        n_Body_y[799] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 800) begin
                        n_Body_x[800] = c_Body_x[799];
                        n_Body_y[800] = c_Body_y[799];
                    end else begin
                        n_Body_x[800] = c_Body_x[c_Size-1];
                        n_Body_y[800] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 801) begin
                        n_Body_x[801] = c_Body_x[800];
                        n_Body_y[801] = c_Body_y[800];
                    end else begin
                        n_Body_x[801] = c_Body_x[c_Size-1];
                        n_Body_y[801] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 802) begin
                        n_Body_x[802] = c_Body_x[801];
                        n_Body_y[802] = c_Body_y[801];
                    end else begin
                        n_Body_x[802] = c_Body_x[c_Size-1];
                        n_Body_y[802] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 803) begin
                        n_Body_x[803] = c_Body_x[802];
                        n_Body_y[803] = c_Body_y[802];
                    end else begin
                        n_Body_x[803] = c_Body_x[c_Size-1];
                        n_Body_y[803] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 804) begin
                        n_Body_x[804] = c_Body_x[803];
                        n_Body_y[804] = c_Body_y[803];
                    end else begin
                        n_Body_x[804] = c_Body_x[c_Size-1];
                        n_Body_y[804] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 805) begin
                        n_Body_x[805] = c_Body_x[804];
                        n_Body_y[805] = c_Body_y[804];
                    end else begin
                        n_Body_x[805] = c_Body_x[c_Size-1];
                        n_Body_y[805] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 806) begin
                        n_Body_x[806] = c_Body_x[805];
                        n_Body_y[806] = c_Body_y[805];
                    end else begin
                        n_Body_x[806] = c_Body_x[c_Size-1];
                        n_Body_y[806] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 807) begin
                        n_Body_x[807] = c_Body_x[806];
                        n_Body_y[807] = c_Body_y[806];
                    end else begin
                        n_Body_x[807] = c_Body_x[c_Size-1];
                        n_Body_y[807] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 808) begin
                        n_Body_x[808] = c_Body_x[807];
                        n_Body_y[808] = c_Body_y[807];
                    end else begin
                        n_Body_x[808] = c_Body_x[c_Size-1];
                        n_Body_y[808] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 809) begin
                        n_Body_x[809] = c_Body_x[808];
                        n_Body_y[809] = c_Body_y[808];
                    end else begin
                        n_Body_x[809] = c_Body_x[c_Size-1];
                        n_Body_y[809] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 810) begin
                        n_Body_x[810] = c_Body_x[809];
                        n_Body_y[810] = c_Body_y[809];
                    end else begin
                        n_Body_x[810] = c_Body_x[c_Size-1];
                        n_Body_y[810] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 811) begin
                        n_Body_x[811] = c_Body_x[810];
                        n_Body_y[811] = c_Body_y[810];
                    end else begin
                        n_Body_x[811] = c_Body_x[c_Size-1];
                        n_Body_y[811] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 812) begin
                        n_Body_x[812] = c_Body_x[811];
                        n_Body_y[812] = c_Body_y[811];
                    end else begin
                        n_Body_x[812] = c_Body_x[c_Size-1];
                        n_Body_y[812] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 813) begin
                        n_Body_x[813] = c_Body_x[812];
                        n_Body_y[813] = c_Body_y[812];
                    end else begin
                        n_Body_x[813] = c_Body_x[c_Size-1];
                        n_Body_y[813] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 814) begin
                        n_Body_x[814] = c_Body_x[813];
                        n_Body_y[814] = c_Body_y[813];
                    end else begin
                        n_Body_x[814] = c_Body_x[c_Size-1];
                        n_Body_y[814] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 815) begin
                        n_Body_x[815] = c_Body_x[814];
                        n_Body_y[815] = c_Body_y[814];
                    end else begin
                        n_Body_x[815] = c_Body_x[c_Size-1];
                        n_Body_y[815] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 816) begin
                        n_Body_x[816] = c_Body_x[815];
                        n_Body_y[816] = c_Body_y[815];
                    end else begin
                        n_Body_x[816] = c_Body_x[c_Size-1];
                        n_Body_y[816] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 817) begin
                        n_Body_x[817] = c_Body_x[816];
                        n_Body_y[817] = c_Body_y[816];
                    end else begin
                        n_Body_x[817] = c_Body_x[c_Size-1];
                        n_Body_y[817] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 818) begin
                        n_Body_x[818] = c_Body_x[817];
                        n_Body_y[818] = c_Body_y[817];
                    end else begin
                        n_Body_x[818] = c_Body_x[c_Size-1];
                        n_Body_y[818] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 819) begin
                        n_Body_x[819] = c_Body_x[818];
                        n_Body_y[819] = c_Body_y[818];
                    end else begin
                        n_Body_x[819] = c_Body_x[c_Size-1];
                        n_Body_y[819] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 820) begin
                        n_Body_x[820] = c_Body_x[819];
                        n_Body_y[820] = c_Body_y[819];
                    end else begin
                        n_Body_x[820] = c_Body_x[c_Size-1];
                        n_Body_y[820] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 821) begin
                        n_Body_x[821] = c_Body_x[820];
                        n_Body_y[821] = c_Body_y[820];
                    end else begin
                        n_Body_x[821] = c_Body_x[c_Size-1];
                        n_Body_y[821] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 822) begin
                        n_Body_x[822] = c_Body_x[821];
                        n_Body_y[822] = c_Body_y[821];
                    end else begin
                        n_Body_x[822] = c_Body_x[c_Size-1];
                        n_Body_y[822] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 823) begin
                        n_Body_x[823] = c_Body_x[822];
                        n_Body_y[823] = c_Body_y[822];
                    end else begin
                        n_Body_x[823] = c_Body_x[c_Size-1];
                        n_Body_y[823] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 824) begin
                        n_Body_x[824] = c_Body_x[823];
                        n_Body_y[824] = c_Body_y[823];
                    end else begin
                        n_Body_x[824] = c_Body_x[c_Size-1];
                        n_Body_y[824] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 825) begin
                        n_Body_x[825] = c_Body_x[824];
                        n_Body_y[825] = c_Body_y[824];
                    end else begin
                        n_Body_x[825] = c_Body_x[c_Size-1];
                        n_Body_y[825] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 826) begin
                        n_Body_x[826] = c_Body_x[825];
                        n_Body_y[826] = c_Body_y[825];
                    end else begin
                        n_Body_x[826] = c_Body_x[c_Size-1];
                        n_Body_y[826] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 827) begin
                        n_Body_x[827] = c_Body_x[826];
                        n_Body_y[827] = c_Body_y[826];
                    end else begin
                        n_Body_x[827] = c_Body_x[c_Size-1];
                        n_Body_y[827] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 828) begin
                        n_Body_x[828] = c_Body_x[827];
                        n_Body_y[828] = c_Body_y[827];
                    end else begin
                        n_Body_x[828] = c_Body_x[c_Size-1];
                        n_Body_y[828] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 829) begin
                        n_Body_x[829] = c_Body_x[828];
                        n_Body_y[829] = c_Body_y[828];
                    end else begin
                        n_Body_x[829] = c_Body_x[c_Size-1];
                        n_Body_y[829] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 830) begin
                        n_Body_x[830] = c_Body_x[829];
                        n_Body_y[830] = c_Body_y[829];
                    end else begin
                        n_Body_x[830] = c_Body_x[c_Size-1];
                        n_Body_y[830] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 831) begin
                        n_Body_x[831] = c_Body_x[830];
                        n_Body_y[831] = c_Body_y[830];
                    end else begin
                        n_Body_x[831] = c_Body_x[c_Size-1];
                        n_Body_y[831] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 832) begin
                        n_Body_x[832] = c_Body_x[831];
                        n_Body_y[832] = c_Body_y[831];
                    end else begin
                        n_Body_x[832] = c_Body_x[c_Size-1];
                        n_Body_y[832] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 833) begin
                        n_Body_x[833] = c_Body_x[832];
                        n_Body_y[833] = c_Body_y[832];
                    end else begin
                        n_Body_x[833] = c_Body_x[c_Size-1];
                        n_Body_y[833] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 834) begin
                        n_Body_x[834] = c_Body_x[833];
                        n_Body_y[834] = c_Body_y[833];
                    end else begin
                        n_Body_x[834] = c_Body_x[c_Size-1];
                        n_Body_y[834] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 835) begin
                        n_Body_x[835] = c_Body_x[834];
                        n_Body_y[835] = c_Body_y[834];
                    end else begin
                        n_Body_x[835] = c_Body_x[c_Size-1];
                        n_Body_y[835] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 836) begin
                        n_Body_x[836] = c_Body_x[835];
                        n_Body_y[836] = c_Body_y[835];
                    end else begin
                        n_Body_x[836] = c_Body_x[c_Size-1];
                        n_Body_y[836] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 837) begin
                        n_Body_x[837] = c_Body_x[836];
                        n_Body_y[837] = c_Body_y[836];
                    end else begin
                        n_Body_x[837] = c_Body_x[c_Size-1];
                        n_Body_y[837] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 838) begin
                        n_Body_x[838] = c_Body_x[837];
                        n_Body_y[838] = c_Body_y[837];
                    end else begin
                        n_Body_x[838] = c_Body_x[c_Size-1];
                        n_Body_y[838] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 839) begin
                        n_Body_x[839] = c_Body_x[838];
                        n_Body_y[839] = c_Body_y[838];
                    end else begin
                        n_Body_x[839] = c_Body_x[c_Size-1];
                        n_Body_y[839] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 840) begin
                        n_Body_x[840] = c_Body_x[839];
                        n_Body_y[840] = c_Body_y[839];
                    end else begin
                        n_Body_x[840] = c_Body_x[c_Size-1];
                        n_Body_y[840] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 841) begin
                        n_Body_x[841] = c_Body_x[840];
                        n_Body_y[841] = c_Body_y[840];
                    end else begin
                        n_Body_x[841] = c_Body_x[c_Size-1];
                        n_Body_y[841] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 842) begin
                        n_Body_x[842] = c_Body_x[841];
                        n_Body_y[842] = c_Body_y[841];
                    end else begin
                        n_Body_x[842] = c_Body_x[c_Size-1];
                        n_Body_y[842] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 843) begin
                        n_Body_x[843] = c_Body_x[842];
                        n_Body_y[843] = c_Body_y[842];
                    end else begin
                        n_Body_x[843] = c_Body_x[c_Size-1];
                        n_Body_y[843] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 844) begin
                        n_Body_x[844] = c_Body_x[843];
                        n_Body_y[844] = c_Body_y[843];
                    end else begin
                        n_Body_x[844] = c_Body_x[c_Size-1];
                        n_Body_y[844] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 845) begin
                        n_Body_x[845] = c_Body_x[844];
                        n_Body_y[845] = c_Body_y[844];
                    end else begin
                        n_Body_x[845] = c_Body_x[c_Size-1];
                        n_Body_y[845] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 846) begin
                        n_Body_x[846] = c_Body_x[845];
                        n_Body_y[846] = c_Body_y[845];
                    end else begin
                        n_Body_x[846] = c_Body_x[c_Size-1];
                        n_Body_y[846] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 847) begin
                        n_Body_x[847] = c_Body_x[846];
                        n_Body_y[847] = c_Body_y[846];
                    end else begin
                        n_Body_x[847] = c_Body_x[c_Size-1];
                        n_Body_y[847] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 848) begin
                        n_Body_x[848] = c_Body_x[847];
                        n_Body_y[848] = c_Body_y[847];
                    end else begin
                        n_Body_x[848] = c_Body_x[c_Size-1];
                        n_Body_y[848] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 849) begin
                        n_Body_x[849] = c_Body_x[848];
                        n_Body_y[849] = c_Body_y[848];
                    end else begin
                        n_Body_x[849] = c_Body_x[c_Size-1];
                        n_Body_y[849] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 850) begin
                        n_Body_x[850] = c_Body_x[849];
                        n_Body_y[850] = c_Body_y[849];
                    end else begin
                        n_Body_x[850] = c_Body_x[c_Size-1];
                        n_Body_y[850] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 851) begin
                        n_Body_x[851] = c_Body_x[850];
                        n_Body_y[851] = c_Body_y[850];
                    end else begin
                        n_Body_x[851] = c_Body_x[c_Size-1];
                        n_Body_y[851] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 852) begin
                        n_Body_x[852] = c_Body_x[851];
                        n_Body_y[852] = c_Body_y[851];
                    end else begin
                        n_Body_x[852] = c_Body_x[c_Size-1];
                        n_Body_y[852] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 853) begin
                        n_Body_x[853] = c_Body_x[852];
                        n_Body_y[853] = c_Body_y[852];
                    end else begin
                        n_Body_x[853] = c_Body_x[c_Size-1];
                        n_Body_y[853] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 854) begin
                        n_Body_x[854] = c_Body_x[853];
                        n_Body_y[854] = c_Body_y[853];
                    end else begin
                        n_Body_x[854] = c_Body_x[c_Size-1];
                        n_Body_y[854] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 855) begin
                        n_Body_x[855] = c_Body_x[854];
                        n_Body_y[855] = c_Body_y[854];
                    end else begin
                        n_Body_x[855] = c_Body_x[c_Size-1];
                        n_Body_y[855] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 856) begin
                        n_Body_x[856] = c_Body_x[855];
                        n_Body_y[856] = c_Body_y[855];
                    end else begin
                        n_Body_x[856] = c_Body_x[c_Size-1];
                        n_Body_y[856] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 857) begin
                        n_Body_x[857] = c_Body_x[856];
                        n_Body_y[857] = c_Body_y[856];
                    end else begin
                        n_Body_x[857] = c_Body_x[c_Size-1];
                        n_Body_y[857] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 858) begin
                        n_Body_x[858] = c_Body_x[857];
                        n_Body_y[858] = c_Body_y[857];
                    end else begin
                        n_Body_x[858] = c_Body_x[c_Size-1];
                        n_Body_y[858] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 859) begin
                        n_Body_x[859] = c_Body_x[858];
                        n_Body_y[859] = c_Body_y[858];
                    end else begin
                        n_Body_x[859] = c_Body_x[c_Size-1];
                        n_Body_y[859] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 860) begin
                        n_Body_x[860] = c_Body_x[859];
                        n_Body_y[860] = c_Body_y[859];
                    end else begin
                        n_Body_x[860] = c_Body_x[c_Size-1];
                        n_Body_y[860] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 861) begin
                        n_Body_x[861] = c_Body_x[860];
                        n_Body_y[861] = c_Body_y[860];
                    end else begin
                        n_Body_x[861] = c_Body_x[c_Size-1];
                        n_Body_y[861] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 862) begin
                        n_Body_x[862] = c_Body_x[861];
                        n_Body_y[862] = c_Body_y[861];
                    end else begin
                        n_Body_x[862] = c_Body_x[c_Size-1];
                        n_Body_y[862] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 863) begin
                        n_Body_x[863] = c_Body_x[862];
                        n_Body_y[863] = c_Body_y[862];
                    end else begin
                        n_Body_x[863] = c_Body_x[c_Size-1];
                        n_Body_y[863] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 864) begin
                        n_Body_x[864] = c_Body_x[863];
                        n_Body_y[864] = c_Body_y[863];
                    end else begin
                        n_Body_x[864] = c_Body_x[c_Size-1];
                        n_Body_y[864] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 865) begin
                        n_Body_x[865] = c_Body_x[864];
                        n_Body_y[865] = c_Body_y[864];
                    end else begin
                        n_Body_x[865] = c_Body_x[c_Size-1];
                        n_Body_y[865] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 866) begin
                        n_Body_x[866] = c_Body_x[865];
                        n_Body_y[866] = c_Body_y[865];
                    end else begin
                        n_Body_x[866] = c_Body_x[c_Size-1];
                        n_Body_y[866] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 867) begin
                        n_Body_x[867] = c_Body_x[866];
                        n_Body_y[867] = c_Body_y[866];
                    end else begin
                        n_Body_x[867] = c_Body_x[c_Size-1];
                        n_Body_y[867] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 868) begin
                        n_Body_x[868] = c_Body_x[867];
                        n_Body_y[868] = c_Body_y[867];
                    end else begin
                        n_Body_x[868] = c_Body_x[c_Size-1];
                        n_Body_y[868] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 869) begin
                        n_Body_x[869] = c_Body_x[868];
                        n_Body_y[869] = c_Body_y[868];
                    end else begin
                        n_Body_x[869] = c_Body_x[c_Size-1];
                        n_Body_y[869] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 870) begin
                        n_Body_x[870] = c_Body_x[869];
                        n_Body_y[870] = c_Body_y[869];
                    end else begin
                        n_Body_x[870] = c_Body_x[c_Size-1];
                        n_Body_y[870] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 871) begin
                        n_Body_x[871] = c_Body_x[870];
                        n_Body_y[871] = c_Body_y[870];
                    end else begin
                        n_Body_x[871] = c_Body_x[c_Size-1];
                        n_Body_y[871] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 872) begin
                        n_Body_x[872] = c_Body_x[871];
                        n_Body_y[872] = c_Body_y[871];
                    end else begin
                        n_Body_x[872] = c_Body_x[c_Size-1];
                        n_Body_y[872] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 873) begin
                        n_Body_x[873] = c_Body_x[872];
                        n_Body_y[873] = c_Body_y[872];
                    end else begin
                        n_Body_x[873] = c_Body_x[c_Size-1];
                        n_Body_y[873] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 874) begin
                        n_Body_x[874] = c_Body_x[873];
                        n_Body_y[874] = c_Body_y[873];
                    end else begin
                        n_Body_x[874] = c_Body_x[c_Size-1];
                        n_Body_y[874] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 875) begin
                        n_Body_x[875] = c_Body_x[874];
                        n_Body_y[875] = c_Body_y[874];
                    end else begin
                        n_Body_x[875] = c_Body_x[c_Size-1];
                        n_Body_y[875] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 876) begin
                        n_Body_x[876] = c_Body_x[875];
                        n_Body_y[876] = c_Body_y[875];
                    end else begin
                        n_Body_x[876] = c_Body_x[c_Size-1];
                        n_Body_y[876] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 877) begin
                        n_Body_x[877] = c_Body_x[876];
                        n_Body_y[877] = c_Body_y[876];
                    end else begin
                        n_Body_x[877] = c_Body_x[c_Size-1];
                        n_Body_y[877] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 878) begin
                        n_Body_x[878] = c_Body_x[877];
                        n_Body_y[878] = c_Body_y[877];
                    end else begin
                        n_Body_x[878] = c_Body_x[c_Size-1];
                        n_Body_y[878] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 879) begin
                        n_Body_x[879] = c_Body_x[878];
                        n_Body_y[879] = c_Body_y[878];
                    end else begin
                        n_Body_x[879] = c_Body_x[c_Size-1];
                        n_Body_y[879] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 880) begin
                        n_Body_x[880] = c_Body_x[879];
                        n_Body_y[880] = c_Body_y[879];
                    end else begin
                        n_Body_x[880] = c_Body_x[c_Size-1];
                        n_Body_y[880] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 881) begin
                        n_Body_x[881] = c_Body_x[880];
                        n_Body_y[881] = c_Body_y[880];
                    end else begin
                        n_Body_x[881] = c_Body_x[c_Size-1];
                        n_Body_y[881] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 882) begin
                        n_Body_x[882] = c_Body_x[881];
                        n_Body_y[882] = c_Body_y[881];
                    end else begin
                        n_Body_x[882] = c_Body_x[c_Size-1];
                        n_Body_y[882] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 883) begin
                        n_Body_x[883] = c_Body_x[882];
                        n_Body_y[883] = c_Body_y[882];
                    end else begin
                        n_Body_x[883] = c_Body_x[c_Size-1];
                        n_Body_y[883] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 884) begin
                        n_Body_x[884] = c_Body_x[883];
                        n_Body_y[884] = c_Body_y[883];
                    end else begin
                        n_Body_x[884] = c_Body_x[c_Size-1];
                        n_Body_y[884] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 885) begin
                        n_Body_x[885] = c_Body_x[884];
                        n_Body_y[885] = c_Body_y[884];
                    end else begin
                        n_Body_x[885] = c_Body_x[c_Size-1];
                        n_Body_y[885] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 886) begin
                        n_Body_x[886] = c_Body_x[885];
                        n_Body_y[886] = c_Body_y[885];
                    end else begin
                        n_Body_x[886] = c_Body_x[c_Size-1];
                        n_Body_y[886] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 887) begin
                        n_Body_x[887] = c_Body_x[886];
                        n_Body_y[887] = c_Body_y[886];
                    end else begin
                        n_Body_x[887] = c_Body_x[c_Size-1];
                        n_Body_y[887] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 888) begin
                        n_Body_x[888] = c_Body_x[887];
                        n_Body_y[888] = c_Body_y[887];
                    end else begin
                        n_Body_x[888] = c_Body_x[c_Size-1];
                        n_Body_y[888] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 889) begin
                        n_Body_x[889] = c_Body_x[888];
                        n_Body_y[889] = c_Body_y[888];
                    end else begin
                        n_Body_x[889] = c_Body_x[c_Size-1];
                        n_Body_y[889] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 890) begin
                        n_Body_x[890] = c_Body_x[889];
                        n_Body_y[890] = c_Body_y[889];
                    end else begin
                        n_Body_x[890] = c_Body_x[c_Size-1];
                        n_Body_y[890] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 891) begin
                        n_Body_x[891] = c_Body_x[890];
                        n_Body_y[891] = c_Body_y[890];
                    end else begin
                        n_Body_x[891] = c_Body_x[c_Size-1];
                        n_Body_y[891] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 892) begin
                        n_Body_x[892] = c_Body_x[891];
                        n_Body_y[892] = c_Body_y[891];
                    end else begin
                        n_Body_x[892] = c_Body_x[c_Size-1];
                        n_Body_y[892] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 893) begin
                        n_Body_x[893] = c_Body_x[892];
                        n_Body_y[893] = c_Body_y[892];
                    end else begin
                        n_Body_x[893] = c_Body_x[c_Size-1];
                        n_Body_y[893] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 894) begin
                        n_Body_x[894] = c_Body_x[893];
                        n_Body_y[894] = c_Body_y[893];
                    end else begin
                        n_Body_x[894] = c_Body_x[c_Size-1];
                        n_Body_y[894] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 895) begin
                        n_Body_x[895] = c_Body_x[894];
                        n_Body_y[895] = c_Body_y[894];
                    end else begin
                        n_Body_x[895] = c_Body_x[c_Size-1];
                        n_Body_y[895] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 896) begin
                        n_Body_x[896] = c_Body_x[895];
                        n_Body_y[896] = c_Body_y[895];
                    end else begin
                        n_Body_x[896] = c_Body_x[c_Size-1];
                        n_Body_y[896] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 897) begin
                        n_Body_x[897] = c_Body_x[896];
                        n_Body_y[897] = c_Body_y[896];
                    end else begin
                        n_Body_x[897] = c_Body_x[c_Size-1];
                        n_Body_y[897] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 898) begin
                        n_Body_x[898] = c_Body_x[897];
                        n_Body_y[898] = c_Body_y[897];
                    end else begin
                        n_Body_x[898] = c_Body_x[c_Size-1];
                        n_Body_y[898] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 899) begin
                        n_Body_x[899] = c_Body_x[898];
                        n_Body_y[899] = c_Body_y[898];
                    end else begin
                        n_Body_x[899] = c_Body_x[c_Size-1];
                        n_Body_y[899] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 900) begin
                        n_Body_x[900] = c_Body_x[899];
                        n_Body_y[900] = c_Body_y[899];
                    end else begin
                        n_Body_x[900] = c_Body_x[c_Size-1];
                        n_Body_y[900] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 901) begin
                        n_Body_x[901] = c_Body_x[900];
                        n_Body_y[901] = c_Body_y[900];
                    end else begin
                        n_Body_x[901] = c_Body_x[c_Size-1];
                        n_Body_y[901] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 902) begin
                        n_Body_x[902] = c_Body_x[901];
                        n_Body_y[902] = c_Body_y[901];
                    end else begin
                        n_Body_x[902] = c_Body_x[c_Size-1];
                        n_Body_y[902] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 903) begin
                        n_Body_x[903] = c_Body_x[902];
                        n_Body_y[903] = c_Body_y[902];
                    end else begin
                        n_Body_x[903] = c_Body_x[c_Size-1];
                        n_Body_y[903] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 904) begin
                        n_Body_x[904] = c_Body_x[903];
                        n_Body_y[904] = c_Body_y[903];
                    end else begin
                        n_Body_x[904] = c_Body_x[c_Size-1];
                        n_Body_y[904] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 905) begin
                        n_Body_x[905] = c_Body_x[904];
                        n_Body_y[905] = c_Body_y[904];
                    end else begin
                        n_Body_x[905] = c_Body_x[c_Size-1];
                        n_Body_y[905] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 906) begin
                        n_Body_x[906] = c_Body_x[905];
                        n_Body_y[906] = c_Body_y[905];
                    end else begin
                        n_Body_x[906] = c_Body_x[c_Size-1];
                        n_Body_y[906] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 907) begin
                        n_Body_x[907] = c_Body_x[906];
                        n_Body_y[907] = c_Body_y[906];
                    end else begin
                        n_Body_x[907] = c_Body_x[c_Size-1];
                        n_Body_y[907] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 908) begin
                        n_Body_x[908] = c_Body_x[907];
                        n_Body_y[908] = c_Body_y[907];
                    end else begin
                        n_Body_x[908] = c_Body_x[c_Size-1];
                        n_Body_y[908] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 909) begin
                        n_Body_x[909] = c_Body_x[908];
                        n_Body_y[909] = c_Body_y[908];
                    end else begin
                        n_Body_x[909] = c_Body_x[c_Size-1];
                        n_Body_y[909] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 910) begin
                        n_Body_x[910] = c_Body_x[909];
                        n_Body_y[910] = c_Body_y[909];
                    end else begin
                        n_Body_x[910] = c_Body_x[c_Size-1];
                        n_Body_y[910] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 911) begin
                        n_Body_x[911] = c_Body_x[910];
                        n_Body_y[911] = c_Body_y[910];
                    end else begin
                        n_Body_x[911] = c_Body_x[c_Size-1];
                        n_Body_y[911] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 912) begin
                        n_Body_x[912] = c_Body_x[911];
                        n_Body_y[912] = c_Body_y[911];
                    end else begin
                        n_Body_x[912] = c_Body_x[c_Size-1];
                        n_Body_y[912] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 913) begin
                        n_Body_x[913] = c_Body_x[912];
                        n_Body_y[913] = c_Body_y[912];
                    end else begin
                        n_Body_x[913] = c_Body_x[c_Size-1];
                        n_Body_y[913] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 914) begin
                        n_Body_x[914] = c_Body_x[913];
                        n_Body_y[914] = c_Body_y[913];
                    end else begin
                        n_Body_x[914] = c_Body_x[c_Size-1];
                        n_Body_y[914] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 915) begin
                        n_Body_x[915] = c_Body_x[914];
                        n_Body_y[915] = c_Body_y[914];
                    end else begin
                        n_Body_x[915] = c_Body_x[c_Size-1];
                        n_Body_y[915] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 916) begin
                        n_Body_x[916] = c_Body_x[915];
                        n_Body_y[916] = c_Body_y[915];
                    end else begin
                        n_Body_x[916] = c_Body_x[c_Size-1];
                        n_Body_y[916] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 917) begin
                        n_Body_x[917] = c_Body_x[916];
                        n_Body_y[917] = c_Body_y[916];
                    end else begin
                        n_Body_x[917] = c_Body_x[c_Size-1];
                        n_Body_y[917] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 918) begin
                        n_Body_x[918] = c_Body_x[917];
                        n_Body_y[918] = c_Body_y[917];
                    end else begin
                        n_Body_x[918] = c_Body_x[c_Size-1];
                        n_Body_y[918] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 919) begin
                        n_Body_x[919] = c_Body_x[918];
                        n_Body_y[919] = c_Body_y[918];
                    end else begin
                        n_Body_x[919] = c_Body_x[c_Size-1];
                        n_Body_y[919] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 920) begin
                        n_Body_x[920] = c_Body_x[919];
                        n_Body_y[920] = c_Body_y[919];
                    end else begin
                        n_Body_x[920] = c_Body_x[c_Size-1];
                        n_Body_y[920] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 921) begin
                        n_Body_x[921] = c_Body_x[920];
                        n_Body_y[921] = c_Body_y[920];
                    end else begin
                        n_Body_x[921] = c_Body_x[c_Size-1];
                        n_Body_y[921] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 922) begin
                        n_Body_x[922] = c_Body_x[921];
                        n_Body_y[922] = c_Body_y[921];
                    end else begin
                        n_Body_x[922] = c_Body_x[c_Size-1];
                        n_Body_y[922] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 923) begin
                        n_Body_x[923] = c_Body_x[922];
                        n_Body_y[923] = c_Body_y[922];
                    end else begin
                        n_Body_x[923] = c_Body_x[c_Size-1];
                        n_Body_y[923] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 924) begin
                        n_Body_x[924] = c_Body_x[923];
                        n_Body_y[924] = c_Body_y[923];
                    end else begin
                        n_Body_x[924] = c_Body_x[c_Size-1];
                        n_Body_y[924] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 925) begin
                        n_Body_x[925] = c_Body_x[924];
                        n_Body_y[925] = c_Body_y[924];
                    end else begin
                        n_Body_x[925] = c_Body_x[c_Size-1];
                        n_Body_y[925] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 926) begin
                        n_Body_x[926] = c_Body_x[925];
                        n_Body_y[926] = c_Body_y[925];
                    end else begin
                        n_Body_x[926] = c_Body_x[c_Size-1];
                        n_Body_y[926] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 927) begin
                        n_Body_x[927] = c_Body_x[926];
                        n_Body_y[927] = c_Body_y[926];
                    end else begin
                        n_Body_x[927] = c_Body_x[c_Size-1];
                        n_Body_y[927] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 928) begin
                        n_Body_x[928] = c_Body_x[927];
                        n_Body_y[928] = c_Body_y[927];
                    end else begin
                        n_Body_x[928] = c_Body_x[c_Size-1];
                        n_Body_y[928] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 929) begin
                        n_Body_x[929] = c_Body_x[928];
                        n_Body_y[929] = c_Body_y[928];
                    end else begin
                        n_Body_x[929] = c_Body_x[c_Size-1];
                        n_Body_y[929] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 930) begin
                        n_Body_x[930] = c_Body_x[929];
                        n_Body_y[930] = c_Body_y[929];
                    end else begin
                        n_Body_x[930] = c_Body_x[c_Size-1];
                        n_Body_y[930] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 931) begin
                        n_Body_x[931] = c_Body_x[930];
                        n_Body_y[931] = c_Body_y[930];
                    end else begin
                        n_Body_x[931] = c_Body_x[c_Size-1];
                        n_Body_y[931] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 932) begin
                        n_Body_x[932] = c_Body_x[931];
                        n_Body_y[932] = c_Body_y[931];
                    end else begin
                        n_Body_x[932] = c_Body_x[c_Size-1];
                        n_Body_y[932] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 933) begin
                        n_Body_x[933] = c_Body_x[932];
                        n_Body_y[933] = c_Body_y[932];
                    end else begin
                        n_Body_x[933] = c_Body_x[c_Size-1];
                        n_Body_y[933] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 934) begin
                        n_Body_x[934] = c_Body_x[933];
                        n_Body_y[934] = c_Body_y[933];
                    end else begin
                        n_Body_x[934] = c_Body_x[c_Size-1];
                        n_Body_y[934] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 935) begin
                        n_Body_x[935] = c_Body_x[934];
                        n_Body_y[935] = c_Body_y[934];
                    end else begin
                        n_Body_x[935] = c_Body_x[c_Size-1];
                        n_Body_y[935] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 936) begin
                        n_Body_x[936] = c_Body_x[935];
                        n_Body_y[936] = c_Body_y[935];
                    end else begin
                        n_Body_x[936] = c_Body_x[c_Size-1];
                        n_Body_y[936] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 937) begin
                        n_Body_x[937] = c_Body_x[936];
                        n_Body_y[937] = c_Body_y[936];
                    end else begin
                        n_Body_x[937] = c_Body_x[c_Size-1];
                        n_Body_y[937] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 938) begin
                        n_Body_x[938] = c_Body_x[937];
                        n_Body_y[938] = c_Body_y[937];
                    end else begin
                        n_Body_x[938] = c_Body_x[c_Size-1];
                        n_Body_y[938] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 939) begin
                        n_Body_x[939] = c_Body_x[938];
                        n_Body_y[939] = c_Body_y[938];
                    end else begin
                        n_Body_x[939] = c_Body_x[c_Size-1];
                        n_Body_y[939] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 940) begin
                        n_Body_x[940] = c_Body_x[939];
                        n_Body_y[940] = c_Body_y[939];
                    end else begin
                        n_Body_x[940] = c_Body_x[c_Size-1];
                        n_Body_y[940] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 941) begin
                        n_Body_x[941] = c_Body_x[940];
                        n_Body_y[941] = c_Body_y[940];
                    end else begin
                        n_Body_x[941] = c_Body_x[c_Size-1];
                        n_Body_y[941] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 942) begin
                        n_Body_x[942] = c_Body_x[941];
                        n_Body_y[942] = c_Body_y[941];
                    end else begin
                        n_Body_x[942] = c_Body_x[c_Size-1];
                        n_Body_y[942] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 943) begin
                        n_Body_x[943] = c_Body_x[942];
                        n_Body_y[943] = c_Body_y[942];
                    end else begin
                        n_Body_x[943] = c_Body_x[c_Size-1];
                        n_Body_y[943] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 944) begin
                        n_Body_x[944] = c_Body_x[943];
                        n_Body_y[944] = c_Body_y[943];
                    end else begin
                        n_Body_x[944] = c_Body_x[c_Size-1];
                        n_Body_y[944] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 945) begin
                        n_Body_x[945] = c_Body_x[944];
                        n_Body_y[945] = c_Body_y[944];
                    end else begin
                        n_Body_x[945] = c_Body_x[c_Size-1];
                        n_Body_y[945] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 946) begin
                        n_Body_x[946] = c_Body_x[945];
                        n_Body_y[946] = c_Body_y[945];
                    end else begin
                        n_Body_x[946] = c_Body_x[c_Size-1];
                        n_Body_y[946] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 947) begin
                        n_Body_x[947] = c_Body_x[946];
                        n_Body_y[947] = c_Body_y[946];
                    end else begin
                        n_Body_x[947] = c_Body_x[c_Size-1];
                        n_Body_y[947] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 948) begin
                        n_Body_x[948] = c_Body_x[947];
                        n_Body_y[948] = c_Body_y[947];
                    end else begin
                        n_Body_x[948] = c_Body_x[c_Size-1];
                        n_Body_y[948] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 949) begin
                        n_Body_x[949] = c_Body_x[948];
                        n_Body_y[949] = c_Body_y[948];
                    end else begin
                        n_Body_x[949] = c_Body_x[c_Size-1];
                        n_Body_y[949] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 950) begin
                        n_Body_x[950] = c_Body_x[949];
                        n_Body_y[950] = c_Body_y[949];
                    end else begin
                        n_Body_x[950] = c_Body_x[c_Size-1];
                        n_Body_y[950] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 951) begin
                        n_Body_x[951] = c_Body_x[950];
                        n_Body_y[951] = c_Body_y[950];
                    end else begin
                        n_Body_x[951] = c_Body_x[c_Size-1];
                        n_Body_y[951] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 952) begin
                        n_Body_x[952] = c_Body_x[951];
                        n_Body_y[952] = c_Body_y[951];
                    end else begin
                        n_Body_x[952] = c_Body_x[c_Size-1];
                        n_Body_y[952] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 953) begin
                        n_Body_x[953] = c_Body_x[952];
                        n_Body_y[953] = c_Body_y[952];
                    end else begin
                        n_Body_x[953] = c_Body_x[c_Size-1];
                        n_Body_y[953] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 954) begin
                        n_Body_x[954] = c_Body_x[953];
                        n_Body_y[954] = c_Body_y[953];
                    end else begin
                        n_Body_x[954] = c_Body_x[c_Size-1];
                        n_Body_y[954] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 955) begin
                        n_Body_x[955] = c_Body_x[954];
                        n_Body_y[955] = c_Body_y[954];
                    end else begin
                        n_Body_x[955] = c_Body_x[c_Size-1];
                        n_Body_y[955] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 956) begin
                        n_Body_x[956] = c_Body_x[955];
                        n_Body_y[956] = c_Body_y[955];
                    end else begin
                        n_Body_x[956] = c_Body_x[c_Size-1];
                        n_Body_y[956] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 957) begin
                        n_Body_x[957] = c_Body_x[956];
                        n_Body_y[957] = c_Body_y[956];
                    end else begin
                        n_Body_x[957] = c_Body_x[c_Size-1];
                        n_Body_y[957] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 958) begin
                        n_Body_x[958] = c_Body_x[957];
                        n_Body_y[958] = c_Body_y[957];
                    end else begin
                        n_Body_x[958] = c_Body_x[c_Size-1];
                        n_Body_y[958] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 959) begin
                        n_Body_x[959] = c_Body_x[958];
                        n_Body_y[959] = c_Body_y[958];
                    end else begin
                        n_Body_x[959] = c_Body_x[c_Size-1];
                        n_Body_y[959] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 960) begin
                        n_Body_x[960] = c_Body_x[959];
                        n_Body_y[960] = c_Body_y[959];
                    end else begin
                        n_Body_x[960] = c_Body_x[c_Size-1];
                        n_Body_y[960] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 961) begin
                        n_Body_x[961] = c_Body_x[960];
                        n_Body_y[961] = c_Body_y[960];
                    end else begin
                        n_Body_x[961] = c_Body_x[c_Size-1];
                        n_Body_y[961] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 962) begin
                        n_Body_x[962] = c_Body_x[961];
                        n_Body_y[962] = c_Body_y[961];
                    end else begin
                        n_Body_x[962] = c_Body_x[c_Size-1];
                        n_Body_y[962] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 963) begin
                        n_Body_x[963] = c_Body_x[962];
                        n_Body_y[963] = c_Body_y[962];
                    end else begin
                        n_Body_x[963] = c_Body_x[c_Size-1];
                        n_Body_y[963] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 964) begin
                        n_Body_x[964] = c_Body_x[963];
                        n_Body_y[964] = c_Body_y[963];
                    end else begin
                        n_Body_x[964] = c_Body_x[c_Size-1];
                        n_Body_y[964] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 965) begin
                        n_Body_x[965] = c_Body_x[964];
                        n_Body_y[965] = c_Body_y[964];
                    end else begin
                        n_Body_x[965] = c_Body_x[c_Size-1];
                        n_Body_y[965] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 966) begin
                        n_Body_x[966] = c_Body_x[965];
                        n_Body_y[966] = c_Body_y[965];
                    end else begin
                        n_Body_x[966] = c_Body_x[c_Size-1];
                        n_Body_y[966] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 967) begin
                        n_Body_x[967] = c_Body_x[966];
                        n_Body_y[967] = c_Body_y[966];
                    end else begin
                        n_Body_x[967] = c_Body_x[c_Size-1];
                        n_Body_y[967] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 968) begin
                        n_Body_x[968] = c_Body_x[967];
                        n_Body_y[968] = c_Body_y[967];
                    end else begin
                        n_Body_x[968] = c_Body_x[c_Size-1];
                        n_Body_y[968] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 969) begin
                        n_Body_x[969] = c_Body_x[968];
                        n_Body_y[969] = c_Body_y[968];
                    end else begin
                        n_Body_x[969] = c_Body_x[c_Size-1];
                        n_Body_y[969] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 970) begin
                        n_Body_x[970] = c_Body_x[969];
                        n_Body_y[970] = c_Body_y[969];
                    end else begin
                        n_Body_x[970] = c_Body_x[c_Size-1];
                        n_Body_y[970] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 971) begin
                        n_Body_x[971] = c_Body_x[970];
                        n_Body_y[971] = c_Body_y[970];
                    end else begin
                        n_Body_x[971] = c_Body_x[c_Size-1];
                        n_Body_y[971] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 972) begin
                        n_Body_x[972] = c_Body_x[971];
                        n_Body_y[972] = c_Body_y[971];
                    end else begin
                        n_Body_x[972] = c_Body_x[c_Size-1];
                        n_Body_y[972] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 973) begin
                        n_Body_x[973] = c_Body_x[972];
                        n_Body_y[973] = c_Body_y[972];
                    end else begin
                        n_Body_x[973] = c_Body_x[c_Size-1];
                        n_Body_y[973] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 974) begin
                        n_Body_x[974] = c_Body_x[973];
                        n_Body_y[974] = c_Body_y[973];
                    end else begin
                        n_Body_x[974] = c_Body_x[c_Size-1];
                        n_Body_y[974] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 975) begin
                        n_Body_x[975] = c_Body_x[974];
                        n_Body_y[975] = c_Body_y[974];
                    end else begin
                        n_Body_x[975] = c_Body_x[c_Size-1];
                        n_Body_y[975] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 976) begin
                        n_Body_x[976] = c_Body_x[975];
                        n_Body_y[976] = c_Body_y[975];
                    end else begin
                        n_Body_x[976] = c_Body_x[c_Size-1];
                        n_Body_y[976] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 977) begin
                        n_Body_x[977] = c_Body_x[976];
                        n_Body_y[977] = c_Body_y[976];
                    end else begin
                        n_Body_x[977] = c_Body_x[c_Size-1];
                        n_Body_y[977] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 978) begin
                        n_Body_x[978] = c_Body_x[977];
                        n_Body_y[978] = c_Body_y[977];
                    end else begin
                        n_Body_x[978] = c_Body_x[c_Size-1];
                        n_Body_y[978] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 979) begin
                        n_Body_x[979] = c_Body_x[978];
                        n_Body_y[979] = c_Body_y[978];
                    end else begin
                        n_Body_x[979] = c_Body_x[c_Size-1];
                        n_Body_y[979] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 980) begin
                        n_Body_x[980] = c_Body_x[979];
                        n_Body_y[980] = c_Body_y[979];
                    end else begin
                        n_Body_x[980] = c_Body_x[c_Size-1];
                        n_Body_y[980] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 981) begin
                        n_Body_x[981] = c_Body_x[980];
                        n_Body_y[981] = c_Body_y[980];
                    end else begin
                        n_Body_x[981] = c_Body_x[c_Size-1];
                        n_Body_y[981] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 982) begin
                        n_Body_x[982] = c_Body_x[981];
                        n_Body_y[982] = c_Body_y[981];
                    end else begin
                        n_Body_x[982] = c_Body_x[c_Size-1];
                        n_Body_y[982] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 983) begin
                        n_Body_x[983] = c_Body_x[982];
                        n_Body_y[983] = c_Body_y[982];
                    end else begin
                        n_Body_x[983] = c_Body_x[c_Size-1];
                        n_Body_y[983] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 984) begin
                        n_Body_x[984] = c_Body_x[983];
                        n_Body_y[984] = c_Body_y[983];
                    end else begin
                        n_Body_x[984] = c_Body_x[c_Size-1];
                        n_Body_y[984] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 985) begin
                        n_Body_x[985] = c_Body_x[984];
                        n_Body_y[985] = c_Body_y[984];
                    end else begin
                        n_Body_x[985] = c_Body_x[c_Size-1];
                        n_Body_y[985] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 986) begin
                        n_Body_x[986] = c_Body_x[985];
                        n_Body_y[986] = c_Body_y[985];
                    end else begin
                        n_Body_x[986] = c_Body_x[c_Size-1];
                        n_Body_y[986] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 987) begin
                        n_Body_x[987] = c_Body_x[986];
                        n_Body_y[987] = c_Body_y[986];
                    end else begin
                        n_Body_x[987] = c_Body_x[c_Size-1];
                        n_Body_y[987] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 988) begin
                        n_Body_x[988] = c_Body_x[987];
                        n_Body_y[988] = c_Body_y[987];
                    end else begin
                        n_Body_x[988] = c_Body_x[c_Size-1];
                        n_Body_y[988] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 989) begin
                        n_Body_x[989] = c_Body_x[988];
                        n_Body_y[989] = c_Body_y[988];
                    end else begin
                        n_Body_x[989] = c_Body_x[c_Size-1];
                        n_Body_y[989] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 990) begin
                        n_Body_x[990] = c_Body_x[989];
                        n_Body_y[990] = c_Body_y[989];
                    end else begin
                        n_Body_x[990] = c_Body_x[c_Size-1];
                        n_Body_y[990] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 991) begin
                        n_Body_x[991] = c_Body_x[990];
                        n_Body_y[991] = c_Body_y[990];
                    end else begin
                        n_Body_x[991] = c_Body_x[c_Size-1];
                        n_Body_y[991] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 992) begin
                        n_Body_x[992] = c_Body_x[991];
                        n_Body_y[992] = c_Body_y[991];
                    end else begin
                        n_Body_x[992] = c_Body_x[c_Size-1];
                        n_Body_y[992] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 993) begin
                        n_Body_x[993] = c_Body_x[992];
                        n_Body_y[993] = c_Body_y[992];
                    end else begin
                        n_Body_x[993] = c_Body_x[c_Size-1];
                        n_Body_y[993] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 994) begin
                        n_Body_x[994] = c_Body_x[993];
                        n_Body_y[994] = c_Body_y[993];
                    end else begin
                        n_Body_x[994] = c_Body_x[c_Size-1];
                        n_Body_y[994] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 995) begin
                        n_Body_x[995] = c_Body_x[994];
                        n_Body_y[995] = c_Body_y[994];
                    end else begin
                        n_Body_x[995] = c_Body_x[c_Size-1];
                        n_Body_y[995] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 996) begin
                        n_Body_x[996] = c_Body_x[995];
                        n_Body_y[996] = c_Body_y[995];
                    end else begin
                        n_Body_x[996] = c_Body_x[c_Size-1];
                        n_Body_y[996] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 997) begin
                        n_Body_x[997] = c_Body_x[996];
                        n_Body_y[997] = c_Body_y[996];
                    end else begin
                        n_Body_x[997] = c_Body_x[c_Size-1];
                        n_Body_y[997] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 998) begin
                        n_Body_x[998] = c_Body_x[997];
                        n_Body_y[998] = c_Body_y[997];
                    end else begin
                        n_Body_x[998] = c_Body_x[c_Size-1];
                        n_Body_y[998] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 999) begin
                        n_Body_x[999] = c_Body_x[998];
                        n_Body_y[999] = c_Body_y[998];
                    end else begin
                        n_Body_x[999] = c_Body_x[c_Size-1];
                        n_Body_y[999] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1000) begin
                        n_Body_x[1000] = c_Body_x[999];
                        n_Body_y[1000] = c_Body_y[999];
                    end else begin
                        n_Body_x[1000] = c_Body_x[c_Size-1];
                        n_Body_y[1000] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1001) begin
                        n_Body_x[1001] = c_Body_x[1000];
                        n_Body_y[1001] = c_Body_y[1000];
                    end else begin
                        n_Body_x[1001] = c_Body_x[c_Size-1];
                        n_Body_y[1001] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1002) begin
                        n_Body_x[1002] = c_Body_x[1001];
                        n_Body_y[1002] = c_Body_y[1001];
                    end else begin
                        n_Body_x[1002] = c_Body_x[c_Size-1];
                        n_Body_y[1002] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1003) begin
                        n_Body_x[1003] = c_Body_x[1002];
                        n_Body_y[1003] = c_Body_y[1002];
                    end else begin
                        n_Body_x[1003] = c_Body_x[c_Size-1];
                        n_Body_y[1003] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1004) begin
                        n_Body_x[1004] = c_Body_x[1003];
                        n_Body_y[1004] = c_Body_y[1003];
                    end else begin
                        n_Body_x[1004] = c_Body_x[c_Size-1];
                        n_Body_y[1004] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1005) begin
                        n_Body_x[1005] = c_Body_x[1004];
                        n_Body_y[1005] = c_Body_y[1004];
                    end else begin
                        n_Body_x[1005] = c_Body_x[c_Size-1];
                        n_Body_y[1005] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1006) begin
                        n_Body_x[1006] = c_Body_x[1005];
                        n_Body_y[1006] = c_Body_y[1005];
                    end else begin
                        n_Body_x[1006] = c_Body_x[c_Size-1];
                        n_Body_y[1006] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1007) begin
                        n_Body_x[1007] = c_Body_x[1006];
                        n_Body_y[1007] = c_Body_y[1006];
                    end else begin
                        n_Body_x[1007] = c_Body_x[c_Size-1];
                        n_Body_y[1007] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1008) begin
                        n_Body_x[1008] = c_Body_x[1007];
                        n_Body_y[1008] = c_Body_y[1007];
                    end else begin
                        n_Body_x[1008] = c_Body_x[c_Size-1];
                        n_Body_y[1008] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1009) begin
                        n_Body_x[1009] = c_Body_x[1008];
                        n_Body_y[1009] = c_Body_y[1008];
                    end else begin
                        n_Body_x[1009] = c_Body_x[c_Size-1];
                        n_Body_y[1009] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1010) begin
                        n_Body_x[1010] = c_Body_x[1009];
                        n_Body_y[1010] = c_Body_y[1009];
                    end else begin
                        n_Body_x[1010] = c_Body_x[c_Size-1];
                        n_Body_y[1010] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1011) begin
                        n_Body_x[1011] = c_Body_x[1010];
                        n_Body_y[1011] = c_Body_y[1010];
                    end else begin
                        n_Body_x[1011] = c_Body_x[c_Size-1];
                        n_Body_y[1011] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1012) begin
                        n_Body_x[1012] = c_Body_x[1011];
                        n_Body_y[1012] = c_Body_y[1011];
                    end else begin
                        n_Body_x[1012] = c_Body_x[c_Size-1];
                        n_Body_y[1012] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1013) begin
                        n_Body_x[1013] = c_Body_x[1012];
                        n_Body_y[1013] = c_Body_y[1012];
                    end else begin
                        n_Body_x[1013] = c_Body_x[c_Size-1];
                        n_Body_y[1013] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1014) begin
                        n_Body_x[1014] = c_Body_x[1013];
                        n_Body_y[1014] = c_Body_y[1013];
                    end else begin
                        n_Body_x[1014] = c_Body_x[c_Size-1];
                        n_Body_y[1014] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1015) begin
                        n_Body_x[1015] = c_Body_x[1014];
                        n_Body_y[1015] = c_Body_y[1014];
                    end else begin
                        n_Body_x[1015] = c_Body_x[c_Size-1];
                        n_Body_y[1015] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1016) begin
                        n_Body_x[1016] = c_Body_x[1015];
                        n_Body_y[1016] = c_Body_y[1015];
                    end else begin
                        n_Body_x[1016] = c_Body_x[c_Size-1];
                        n_Body_y[1016] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1017) begin
                        n_Body_x[1017] = c_Body_x[1016];
                        n_Body_y[1017] = c_Body_y[1016];
                    end else begin
                        n_Body_x[1017] = c_Body_x[c_Size-1];
                        n_Body_y[1017] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1018) begin
                        n_Body_x[1018] = c_Body_x[1017];
                        n_Body_y[1018] = c_Body_y[1017];
                    end else begin
                        n_Body_x[1018] = c_Body_x[c_Size-1];
                        n_Body_y[1018] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1019) begin
                        n_Body_x[1019] = c_Body_x[1018];
                        n_Body_y[1019] = c_Body_y[1018];
                    end else begin
                        n_Body_x[1019] = c_Body_x[c_Size-1];
                        n_Body_y[1019] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1020) begin
                        n_Body_x[1020] = c_Body_x[1019];
                        n_Body_y[1020] = c_Body_y[1019];
                    end else begin
                        n_Body_x[1020] = c_Body_x[c_Size-1];
                        n_Body_y[1020] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1021) begin
                        n_Body_x[1021] = c_Body_x[1020];
                        n_Body_y[1021] = c_Body_y[1020];
                    end else begin
                        n_Body_x[1021] = c_Body_x[c_Size-1];
                        n_Body_y[1021] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1022) begin
                        n_Body_x[1022] = c_Body_x[1021];
                        n_Body_y[1022] = c_Body_y[1021];
                    end else begin
                        n_Body_x[1022] = c_Body_x[c_Size-1];
                        n_Body_y[1022] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1023) begin
                        n_Body_x[1023] = c_Body_x[1022];
                        n_Body_y[1023] = c_Body_y[1022];
                    end else begin
                        n_Body_x[1023] = c_Body_x[c_Size-1];
                        n_Body_y[1023] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1024) begin
                        n_Body_x[1024] = c_Body_x[1023];
                        n_Body_y[1024] = c_Body_y[1023];
                    end else begin
                        n_Body_x[1024] = c_Body_x[c_Size-1];
                        n_Body_y[1024] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1025) begin
                        n_Body_x[1025] = c_Body_x[1024];
                        n_Body_y[1025] = c_Body_y[1024];
                    end else begin
                        n_Body_x[1025] = c_Body_x[c_Size-1];
                        n_Body_y[1025] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1026) begin
                        n_Body_x[1026] = c_Body_x[1025];
                        n_Body_y[1026] = c_Body_y[1025];
                    end else begin
                        n_Body_x[1026] = c_Body_x[c_Size-1];
                        n_Body_y[1026] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1027) begin
                        n_Body_x[1027] = c_Body_x[1026];
                        n_Body_y[1027] = c_Body_y[1026];
                    end else begin
                        n_Body_x[1027] = c_Body_x[c_Size-1];
                        n_Body_y[1027] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1028) begin
                        n_Body_x[1028] = c_Body_x[1027];
                        n_Body_y[1028] = c_Body_y[1027];
                    end else begin
                        n_Body_x[1028] = c_Body_x[c_Size-1];
                        n_Body_y[1028] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1029) begin
                        n_Body_x[1029] = c_Body_x[1028];
                        n_Body_y[1029] = c_Body_y[1028];
                    end else begin
                        n_Body_x[1029] = c_Body_x[c_Size-1];
                        n_Body_y[1029] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1030) begin
                        n_Body_x[1030] = c_Body_x[1029];
                        n_Body_y[1030] = c_Body_y[1029];
                    end else begin
                        n_Body_x[1030] = c_Body_x[c_Size-1];
                        n_Body_y[1030] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1031) begin
                        n_Body_x[1031] = c_Body_x[1030];
                        n_Body_y[1031] = c_Body_y[1030];
                    end else begin
                        n_Body_x[1031] = c_Body_x[c_Size-1];
                        n_Body_y[1031] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1032) begin
                        n_Body_x[1032] = c_Body_x[1031];
                        n_Body_y[1032] = c_Body_y[1031];
                    end else begin
                        n_Body_x[1032] = c_Body_x[c_Size-1];
                        n_Body_y[1032] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1033) begin
                        n_Body_x[1033] = c_Body_x[1032];
                        n_Body_y[1033] = c_Body_y[1032];
                    end else begin
                        n_Body_x[1033] = c_Body_x[c_Size-1];
                        n_Body_y[1033] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1034) begin
                        n_Body_x[1034] = c_Body_x[1033];
                        n_Body_y[1034] = c_Body_y[1033];
                    end else begin
                        n_Body_x[1034] = c_Body_x[c_Size-1];
                        n_Body_y[1034] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1035) begin
                        n_Body_x[1035] = c_Body_x[1034];
                        n_Body_y[1035] = c_Body_y[1034];
                    end else begin
                        n_Body_x[1035] = c_Body_x[c_Size-1];
                        n_Body_y[1035] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1036) begin
                        n_Body_x[1036] = c_Body_x[1035];
                        n_Body_y[1036] = c_Body_y[1035];
                    end else begin
                        n_Body_x[1036] = c_Body_x[c_Size-1];
                        n_Body_y[1036] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1037) begin
                        n_Body_x[1037] = c_Body_x[1036];
                        n_Body_y[1037] = c_Body_y[1036];
                    end else begin
                        n_Body_x[1037] = c_Body_x[c_Size-1];
                        n_Body_y[1037] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1038) begin
                        n_Body_x[1038] = c_Body_x[1037];
                        n_Body_y[1038] = c_Body_y[1037];
                    end else begin
                        n_Body_x[1038] = c_Body_x[c_Size-1];
                        n_Body_y[1038] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1039) begin
                        n_Body_x[1039] = c_Body_x[1038];
                        n_Body_y[1039] = c_Body_y[1038];
                    end else begin
                        n_Body_x[1039] = c_Body_x[c_Size-1];
                        n_Body_y[1039] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1040) begin
                        n_Body_x[1040] = c_Body_x[1039];
                        n_Body_y[1040] = c_Body_y[1039];
                    end else begin
                        n_Body_x[1040] = c_Body_x[c_Size-1];
                        n_Body_y[1040] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1041) begin
                        n_Body_x[1041] = c_Body_x[1040];
                        n_Body_y[1041] = c_Body_y[1040];
                    end else begin
                        n_Body_x[1041] = c_Body_x[c_Size-1];
                        n_Body_y[1041] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1042) begin
                        n_Body_x[1042] = c_Body_x[1041];
                        n_Body_y[1042] = c_Body_y[1041];
                    end else begin
                        n_Body_x[1042] = c_Body_x[c_Size-1];
                        n_Body_y[1042] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1043) begin
                        n_Body_x[1043] = c_Body_x[1042];
                        n_Body_y[1043] = c_Body_y[1042];
                    end else begin
                        n_Body_x[1043] = c_Body_x[c_Size-1];
                        n_Body_y[1043] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1044) begin
                        n_Body_x[1044] = c_Body_x[1043];
                        n_Body_y[1044] = c_Body_y[1043];
                    end else begin
                        n_Body_x[1044] = c_Body_x[c_Size-1];
                        n_Body_y[1044] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1045) begin
                        n_Body_x[1045] = c_Body_x[1044];
                        n_Body_y[1045] = c_Body_y[1044];
                    end else begin
                        n_Body_x[1045] = c_Body_x[c_Size-1];
                        n_Body_y[1045] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1046) begin
                        n_Body_x[1046] = c_Body_x[1045];
                        n_Body_y[1046] = c_Body_y[1045];
                    end else begin
                        n_Body_x[1046] = c_Body_x[c_Size-1];
                        n_Body_y[1046] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1047) begin
                        n_Body_x[1047] = c_Body_x[1046];
                        n_Body_y[1047] = c_Body_y[1046];
                    end else begin
                        n_Body_x[1047] = c_Body_x[c_Size-1];
                        n_Body_y[1047] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1048) begin
                        n_Body_x[1048] = c_Body_x[1047];
                        n_Body_y[1048] = c_Body_y[1047];
                    end else begin
                        n_Body_x[1048] = c_Body_x[c_Size-1];
                        n_Body_y[1048] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1049) begin
                        n_Body_x[1049] = c_Body_x[1048];
                        n_Body_y[1049] = c_Body_y[1048];
                    end else begin
                        n_Body_x[1049] = c_Body_x[c_Size-1];
                        n_Body_y[1049] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1050) begin
                        n_Body_x[1050] = c_Body_x[1049];
                        n_Body_y[1050] = c_Body_y[1049];
                    end else begin
                        n_Body_x[1050] = c_Body_x[c_Size-1];
                        n_Body_y[1050] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1051) begin
                        n_Body_x[1051] = c_Body_x[1050];
                        n_Body_y[1051] = c_Body_y[1050];
                    end else begin
                        n_Body_x[1051] = c_Body_x[c_Size-1];
                        n_Body_y[1051] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1052) begin
                        n_Body_x[1052] = c_Body_x[1051];
                        n_Body_y[1052] = c_Body_y[1051];
                    end else begin
                        n_Body_x[1052] = c_Body_x[c_Size-1];
                        n_Body_y[1052] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1053) begin
                        n_Body_x[1053] = c_Body_x[1052];
                        n_Body_y[1053] = c_Body_y[1052];
                    end else begin
                        n_Body_x[1053] = c_Body_x[c_Size-1];
                        n_Body_y[1053] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1054) begin
                        n_Body_x[1054] = c_Body_x[1053];
                        n_Body_y[1054] = c_Body_y[1053];
                    end else begin
                        n_Body_x[1054] = c_Body_x[c_Size-1];
                        n_Body_y[1054] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1055) begin
                        n_Body_x[1055] = c_Body_x[1054];
                        n_Body_y[1055] = c_Body_y[1054];
                    end else begin
                        n_Body_x[1055] = c_Body_x[c_Size-1];
                        n_Body_y[1055] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1056) begin
                        n_Body_x[1056] = c_Body_x[1055];
                        n_Body_y[1056] = c_Body_y[1055];
                    end else begin
                        n_Body_x[1056] = c_Body_x[c_Size-1];
                        n_Body_y[1056] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1057) begin
                        n_Body_x[1057] = c_Body_x[1056];
                        n_Body_y[1057] = c_Body_y[1056];
                    end else begin
                        n_Body_x[1057] = c_Body_x[c_Size-1];
                        n_Body_y[1057] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1058) begin
                        n_Body_x[1058] = c_Body_x[1057];
                        n_Body_y[1058] = c_Body_y[1057];
                    end else begin
                        n_Body_x[1058] = c_Body_x[c_Size-1];
                        n_Body_y[1058] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1059) begin
                        n_Body_x[1059] = c_Body_x[1058];
                        n_Body_y[1059] = c_Body_y[1058];
                    end else begin
                        n_Body_x[1059] = c_Body_x[c_Size-1];
                        n_Body_y[1059] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1060) begin
                        n_Body_x[1060] = c_Body_x[1059];
                        n_Body_y[1060] = c_Body_y[1059];
                    end else begin
                        n_Body_x[1060] = c_Body_x[c_Size-1];
                        n_Body_y[1060] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1061) begin
                        n_Body_x[1061] = c_Body_x[1060];
                        n_Body_y[1061] = c_Body_y[1060];
                    end else begin
                        n_Body_x[1061] = c_Body_x[c_Size-1];
                        n_Body_y[1061] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1062) begin
                        n_Body_x[1062] = c_Body_x[1061];
                        n_Body_y[1062] = c_Body_y[1061];
                    end else begin
                        n_Body_x[1062] = c_Body_x[c_Size-1];
                        n_Body_y[1062] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1063) begin
                        n_Body_x[1063] = c_Body_x[1062];
                        n_Body_y[1063] = c_Body_y[1062];
                    end else begin
                        n_Body_x[1063] = c_Body_x[c_Size-1];
                        n_Body_y[1063] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1064) begin
                        n_Body_x[1064] = c_Body_x[1063];
                        n_Body_y[1064] = c_Body_y[1063];
                    end else begin
                        n_Body_x[1064] = c_Body_x[c_Size-1];
                        n_Body_y[1064] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1065) begin
                        n_Body_x[1065] = c_Body_x[1064];
                        n_Body_y[1065] = c_Body_y[1064];
                    end else begin
                        n_Body_x[1065] = c_Body_x[c_Size-1];
                        n_Body_y[1065] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1066) begin
                        n_Body_x[1066] = c_Body_x[1065];
                        n_Body_y[1066] = c_Body_y[1065];
                    end else begin
                        n_Body_x[1066] = c_Body_x[c_Size-1];
                        n_Body_y[1066] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1067) begin
                        n_Body_x[1067] = c_Body_x[1066];
                        n_Body_y[1067] = c_Body_y[1066];
                    end else begin
                        n_Body_x[1067] = c_Body_x[c_Size-1];
                        n_Body_y[1067] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1068) begin
                        n_Body_x[1068] = c_Body_x[1067];
                        n_Body_y[1068] = c_Body_y[1067];
                    end else begin
                        n_Body_x[1068] = c_Body_x[c_Size-1];
                        n_Body_y[1068] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1069) begin
                        n_Body_x[1069] = c_Body_x[1068];
                        n_Body_y[1069] = c_Body_y[1068];
                    end else begin
                        n_Body_x[1069] = c_Body_x[c_Size-1];
                        n_Body_y[1069] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1070) begin
                        n_Body_x[1070] = c_Body_x[1069];
                        n_Body_y[1070] = c_Body_y[1069];
                    end else begin
                        n_Body_x[1070] = c_Body_x[c_Size-1];
                        n_Body_y[1070] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1071) begin
                        n_Body_x[1071] = c_Body_x[1070];
                        n_Body_y[1071] = c_Body_y[1070];
                    end else begin
                        n_Body_x[1071] = c_Body_x[c_Size-1];
                        n_Body_y[1071] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1072) begin
                        n_Body_x[1072] = c_Body_x[1071];
                        n_Body_y[1072] = c_Body_y[1071];
                    end else begin
                        n_Body_x[1072] = c_Body_x[c_Size-1];
                        n_Body_y[1072] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1073) begin
                        n_Body_x[1073] = c_Body_x[1072];
                        n_Body_y[1073] = c_Body_y[1072];
                    end else begin
                        n_Body_x[1073] = c_Body_x[c_Size-1];
                        n_Body_y[1073] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1074) begin
                        n_Body_x[1074] = c_Body_x[1073];
                        n_Body_y[1074] = c_Body_y[1073];
                    end else begin
                        n_Body_x[1074] = c_Body_x[c_Size-1];
                        n_Body_y[1074] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1075) begin
                        n_Body_x[1075] = c_Body_x[1074];
                        n_Body_y[1075] = c_Body_y[1074];
                    end else begin
                        n_Body_x[1075] = c_Body_x[c_Size-1];
                        n_Body_y[1075] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1076) begin
                        n_Body_x[1076] = c_Body_x[1075];
                        n_Body_y[1076] = c_Body_y[1075];
                    end else begin
                        n_Body_x[1076] = c_Body_x[c_Size-1];
                        n_Body_y[1076] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1077) begin
                        n_Body_x[1077] = c_Body_x[1076];
                        n_Body_y[1077] = c_Body_y[1076];
                    end else begin
                        n_Body_x[1077] = c_Body_x[c_Size-1];
                        n_Body_y[1077] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1078) begin
                        n_Body_x[1078] = c_Body_x[1077];
                        n_Body_y[1078] = c_Body_y[1077];
                    end else begin
                        n_Body_x[1078] = c_Body_x[c_Size-1];
                        n_Body_y[1078] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1079) begin
                        n_Body_x[1079] = c_Body_x[1078];
                        n_Body_y[1079] = c_Body_y[1078];
                    end else begin
                        n_Body_x[1079] = c_Body_x[c_Size-1];
                        n_Body_y[1079] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1080) begin
                        n_Body_x[1080] = c_Body_x[1079];
                        n_Body_y[1080] = c_Body_y[1079];
                    end else begin
                        n_Body_x[1080] = c_Body_x[c_Size-1];
                        n_Body_y[1080] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1081) begin
                        n_Body_x[1081] = c_Body_x[1080];
                        n_Body_y[1081] = c_Body_y[1080];
                    end else begin
                        n_Body_x[1081] = c_Body_x[c_Size-1];
                        n_Body_y[1081] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1082) begin
                        n_Body_x[1082] = c_Body_x[1081];
                        n_Body_y[1082] = c_Body_y[1081];
                    end else begin
                        n_Body_x[1082] = c_Body_x[c_Size-1];
                        n_Body_y[1082] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1083) begin
                        n_Body_x[1083] = c_Body_x[1082];
                        n_Body_y[1083] = c_Body_y[1082];
                    end else begin
                        n_Body_x[1083] = c_Body_x[c_Size-1];
                        n_Body_y[1083] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1084) begin
                        n_Body_x[1084] = c_Body_x[1083];
                        n_Body_y[1084] = c_Body_y[1083];
                    end else begin
                        n_Body_x[1084] = c_Body_x[c_Size-1];
                        n_Body_y[1084] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1085) begin
                        n_Body_x[1085] = c_Body_x[1084];
                        n_Body_y[1085] = c_Body_y[1084];
                    end else begin
                        n_Body_x[1085] = c_Body_x[c_Size-1];
                        n_Body_y[1085] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1086) begin
                        n_Body_x[1086] = c_Body_x[1085];
                        n_Body_y[1086] = c_Body_y[1085];
                    end else begin
                        n_Body_x[1086] = c_Body_x[c_Size-1];
                        n_Body_y[1086] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1087) begin
                        n_Body_x[1087] = c_Body_x[1086];
                        n_Body_y[1087] = c_Body_y[1086];
                    end else begin
                        n_Body_x[1087] = c_Body_x[c_Size-1];
                        n_Body_y[1087] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1088) begin
                        n_Body_x[1088] = c_Body_x[1087];
                        n_Body_y[1088] = c_Body_y[1087];
                    end else begin
                        n_Body_x[1088] = c_Body_x[c_Size-1];
                        n_Body_y[1088] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1089) begin
                        n_Body_x[1089] = c_Body_x[1088];
                        n_Body_y[1089] = c_Body_y[1088];
                    end else begin
                        n_Body_x[1089] = c_Body_x[c_Size-1];
                        n_Body_y[1089] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1090) begin
                        n_Body_x[1090] = c_Body_x[1089];
                        n_Body_y[1090] = c_Body_y[1089];
                    end else begin
                        n_Body_x[1090] = c_Body_x[c_Size-1];
                        n_Body_y[1090] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1091) begin
                        n_Body_x[1091] = c_Body_x[1090];
                        n_Body_y[1091] = c_Body_y[1090];
                    end else begin
                        n_Body_x[1091] = c_Body_x[c_Size-1];
                        n_Body_y[1091] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1092) begin
                        n_Body_x[1092] = c_Body_x[1091];
                        n_Body_y[1092] = c_Body_y[1091];
                    end else begin
                        n_Body_x[1092] = c_Body_x[c_Size-1];
                        n_Body_y[1092] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1093) begin
                        n_Body_x[1093] = c_Body_x[1092];
                        n_Body_y[1093] = c_Body_y[1092];
                    end else begin
                        n_Body_x[1093] = c_Body_x[c_Size-1];
                        n_Body_y[1093] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1094) begin
                        n_Body_x[1094] = c_Body_x[1093];
                        n_Body_y[1094] = c_Body_y[1093];
                    end else begin
                        n_Body_x[1094] = c_Body_x[c_Size-1];
                        n_Body_y[1094] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1095) begin
                        n_Body_x[1095] = c_Body_x[1094];
                        n_Body_y[1095] = c_Body_y[1094];
                    end else begin
                        n_Body_x[1095] = c_Body_x[c_Size-1];
                        n_Body_y[1095] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1096) begin
                        n_Body_x[1096] = c_Body_x[1095];
                        n_Body_y[1096] = c_Body_y[1095];
                    end else begin
                        n_Body_x[1096] = c_Body_x[c_Size-1];
                        n_Body_y[1096] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1097) begin
                        n_Body_x[1097] = c_Body_x[1096];
                        n_Body_y[1097] = c_Body_y[1096];
                    end else begin
                        n_Body_x[1097] = c_Body_x[c_Size-1];
                        n_Body_y[1097] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1098) begin
                        n_Body_x[1098] = c_Body_x[1097];
                        n_Body_y[1098] = c_Body_y[1097];
                    end else begin
                        n_Body_x[1098] = c_Body_x[c_Size-1];
                        n_Body_y[1098] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1099) begin
                        n_Body_x[1099] = c_Body_x[1098];
                        n_Body_y[1099] = c_Body_y[1098];
                    end else begin
                        n_Body_x[1099] = c_Body_x[c_Size-1];
                        n_Body_y[1099] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1100) begin
                        n_Body_x[1100] = c_Body_x[1099];
                        n_Body_y[1100] = c_Body_y[1099];
                    end else begin
                        n_Body_x[1100] = c_Body_x[c_Size-1];
                        n_Body_y[1100] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1101) begin
                        n_Body_x[1101] = c_Body_x[1100];
                        n_Body_y[1101] = c_Body_y[1100];
                    end else begin
                        n_Body_x[1101] = c_Body_x[c_Size-1];
                        n_Body_y[1101] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1102) begin
                        n_Body_x[1102] = c_Body_x[1101];
                        n_Body_y[1102] = c_Body_y[1101];
                    end else begin
                        n_Body_x[1102] = c_Body_x[c_Size-1];
                        n_Body_y[1102] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1103) begin
                        n_Body_x[1103] = c_Body_x[1102];
                        n_Body_y[1103] = c_Body_y[1102];
                    end else begin
                        n_Body_x[1103] = c_Body_x[c_Size-1];
                        n_Body_y[1103] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1104) begin
                        n_Body_x[1104] = c_Body_x[1103];
                        n_Body_y[1104] = c_Body_y[1103];
                    end else begin
                        n_Body_x[1104] = c_Body_x[c_Size-1];
                        n_Body_y[1104] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1105) begin
                        n_Body_x[1105] = c_Body_x[1104];
                        n_Body_y[1105] = c_Body_y[1104];
                    end else begin
                        n_Body_x[1105] = c_Body_x[c_Size-1];
                        n_Body_y[1105] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1106) begin
                        n_Body_x[1106] = c_Body_x[1105];
                        n_Body_y[1106] = c_Body_y[1105];
                    end else begin
                        n_Body_x[1106] = c_Body_x[c_Size-1];
                        n_Body_y[1106] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1107) begin
                        n_Body_x[1107] = c_Body_x[1106];
                        n_Body_y[1107] = c_Body_y[1106];
                    end else begin
                        n_Body_x[1107] = c_Body_x[c_Size-1];
                        n_Body_y[1107] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1108) begin
                        n_Body_x[1108] = c_Body_x[1107];
                        n_Body_y[1108] = c_Body_y[1107];
                    end else begin
                        n_Body_x[1108] = c_Body_x[c_Size-1];
                        n_Body_y[1108] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1109) begin
                        n_Body_x[1109] = c_Body_x[1108];
                        n_Body_y[1109] = c_Body_y[1108];
                    end else begin
                        n_Body_x[1109] = c_Body_x[c_Size-1];
                        n_Body_y[1109] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1110) begin
                        n_Body_x[1110] = c_Body_x[1109];
                        n_Body_y[1110] = c_Body_y[1109];
                    end else begin
                        n_Body_x[1110] = c_Body_x[c_Size-1];
                        n_Body_y[1110] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1111) begin
                        n_Body_x[1111] = c_Body_x[1110];
                        n_Body_y[1111] = c_Body_y[1110];
                    end else begin
                        n_Body_x[1111] = c_Body_x[c_Size-1];
                        n_Body_y[1111] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1112) begin
                        n_Body_x[1112] = c_Body_x[1111];
                        n_Body_y[1112] = c_Body_y[1111];
                    end else begin
                        n_Body_x[1112] = c_Body_x[c_Size-1];
                        n_Body_y[1112] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1113) begin
                        n_Body_x[1113] = c_Body_x[1112];
                        n_Body_y[1113] = c_Body_y[1112];
                    end else begin
                        n_Body_x[1113] = c_Body_x[c_Size-1];
                        n_Body_y[1113] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1114) begin
                        n_Body_x[1114] = c_Body_x[1113];
                        n_Body_y[1114] = c_Body_y[1113];
                    end else begin
                        n_Body_x[1114] = c_Body_x[c_Size-1];
                        n_Body_y[1114] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1115) begin
                        n_Body_x[1115] = c_Body_x[1114];
                        n_Body_y[1115] = c_Body_y[1114];
                    end else begin
                        n_Body_x[1115] = c_Body_x[c_Size-1];
                        n_Body_y[1115] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1116) begin
                        n_Body_x[1116] = c_Body_x[1115];
                        n_Body_y[1116] = c_Body_y[1115];
                    end else begin
                        n_Body_x[1116] = c_Body_x[c_Size-1];
                        n_Body_y[1116] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1117) begin
                        n_Body_x[1117] = c_Body_x[1116];
                        n_Body_y[1117] = c_Body_y[1116];
                    end else begin
                        n_Body_x[1117] = c_Body_x[c_Size-1];
                        n_Body_y[1117] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1118) begin
                        n_Body_x[1118] = c_Body_x[1117];
                        n_Body_y[1118] = c_Body_y[1117];
                    end else begin
                        n_Body_x[1118] = c_Body_x[c_Size-1];
                        n_Body_y[1118] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1119) begin
                        n_Body_x[1119] = c_Body_x[1118];
                        n_Body_y[1119] = c_Body_y[1118];
                    end else begin
                        n_Body_x[1119] = c_Body_x[c_Size-1];
                        n_Body_y[1119] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1120) begin
                        n_Body_x[1120] = c_Body_x[1119];
                        n_Body_y[1120] = c_Body_y[1119];
                    end else begin
                        n_Body_x[1120] = c_Body_x[c_Size-1];
                        n_Body_y[1120] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1121) begin
                        n_Body_x[1121] = c_Body_x[1120];
                        n_Body_y[1121] = c_Body_y[1120];
                    end else begin
                        n_Body_x[1121] = c_Body_x[c_Size-1];
                        n_Body_y[1121] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1122) begin
                        n_Body_x[1122] = c_Body_x[1121];
                        n_Body_y[1122] = c_Body_y[1121];
                    end else begin
                        n_Body_x[1122] = c_Body_x[c_Size-1];
                        n_Body_y[1122] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1123) begin
                        n_Body_x[1123] = c_Body_x[1122];
                        n_Body_y[1123] = c_Body_y[1122];
                    end else begin
                        n_Body_x[1123] = c_Body_x[c_Size-1];
                        n_Body_y[1123] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1124) begin
                        n_Body_x[1124] = c_Body_x[1123];
                        n_Body_y[1124] = c_Body_y[1123];
                    end else begin
                        n_Body_x[1124] = c_Body_x[c_Size-1];
                        n_Body_y[1124] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1125) begin
                        n_Body_x[1125] = c_Body_x[1124];
                        n_Body_y[1125] = c_Body_y[1124];
                    end else begin
                        n_Body_x[1125] = c_Body_x[c_Size-1];
                        n_Body_y[1125] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1126) begin
                        n_Body_x[1126] = c_Body_x[1125];
                        n_Body_y[1126] = c_Body_y[1125];
                    end else begin
                        n_Body_x[1126] = c_Body_x[c_Size-1];
                        n_Body_y[1126] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1127) begin
                        n_Body_x[1127] = c_Body_x[1126];
                        n_Body_y[1127] = c_Body_y[1126];
                    end else begin
                        n_Body_x[1127] = c_Body_x[c_Size-1];
                        n_Body_y[1127] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1128) begin
                        n_Body_x[1128] = c_Body_x[1127];
                        n_Body_y[1128] = c_Body_y[1127];
                    end else begin
                        n_Body_x[1128] = c_Body_x[c_Size-1];
                        n_Body_y[1128] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1129) begin
                        n_Body_x[1129] = c_Body_x[1128];
                        n_Body_y[1129] = c_Body_y[1128];
                    end else begin
                        n_Body_x[1129] = c_Body_x[c_Size-1];
                        n_Body_y[1129] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1130) begin
                        n_Body_x[1130] = c_Body_x[1129];
                        n_Body_y[1130] = c_Body_y[1129];
                    end else begin
                        n_Body_x[1130] = c_Body_x[c_Size-1];
                        n_Body_y[1130] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1131) begin
                        n_Body_x[1131] = c_Body_x[1130];
                        n_Body_y[1131] = c_Body_y[1130];
                    end else begin
                        n_Body_x[1131] = c_Body_x[c_Size-1];
                        n_Body_y[1131] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1132) begin
                        n_Body_x[1132] = c_Body_x[1131];
                        n_Body_y[1132] = c_Body_y[1131];
                    end else begin
                        n_Body_x[1132] = c_Body_x[c_Size-1];
                        n_Body_y[1132] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1133) begin
                        n_Body_x[1133] = c_Body_x[1132];
                        n_Body_y[1133] = c_Body_y[1132];
                    end else begin
                        n_Body_x[1133] = c_Body_x[c_Size-1];
                        n_Body_y[1133] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1134) begin
                        n_Body_x[1134] = c_Body_x[1133];
                        n_Body_y[1134] = c_Body_y[1133];
                    end else begin
                        n_Body_x[1134] = c_Body_x[c_Size-1];
                        n_Body_y[1134] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1135) begin
                        n_Body_x[1135] = c_Body_x[1134];
                        n_Body_y[1135] = c_Body_y[1134];
                    end else begin
                        n_Body_x[1135] = c_Body_x[c_Size-1];
                        n_Body_y[1135] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1136) begin
                        n_Body_x[1136] = c_Body_x[1135];
                        n_Body_y[1136] = c_Body_y[1135];
                    end else begin
                        n_Body_x[1136] = c_Body_x[c_Size-1];
                        n_Body_y[1136] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1137) begin
                        n_Body_x[1137] = c_Body_x[1136];
                        n_Body_y[1137] = c_Body_y[1136];
                    end else begin
                        n_Body_x[1137] = c_Body_x[c_Size-1];
                        n_Body_y[1137] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1138) begin
                        n_Body_x[1138] = c_Body_x[1137];
                        n_Body_y[1138] = c_Body_y[1137];
                    end else begin
                        n_Body_x[1138] = c_Body_x[c_Size-1];
                        n_Body_y[1138] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1139) begin
                        n_Body_x[1139] = c_Body_x[1138];
                        n_Body_y[1139] = c_Body_y[1138];
                    end else begin
                        n_Body_x[1139] = c_Body_x[c_Size-1];
                        n_Body_y[1139] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1140) begin
                        n_Body_x[1140] = c_Body_x[1139];
                        n_Body_y[1140] = c_Body_y[1139];
                    end else begin
                        n_Body_x[1140] = c_Body_x[c_Size-1];
                        n_Body_y[1140] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1141) begin
                        n_Body_x[1141] = c_Body_x[1140];
                        n_Body_y[1141] = c_Body_y[1140];
                    end else begin
                        n_Body_x[1141] = c_Body_x[c_Size-1];
                        n_Body_y[1141] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1142) begin
                        n_Body_x[1142] = c_Body_x[1141];
                        n_Body_y[1142] = c_Body_y[1141];
                    end else begin
                        n_Body_x[1142] = c_Body_x[c_Size-1];
                        n_Body_y[1142] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1143) begin
                        n_Body_x[1143] = c_Body_x[1142];
                        n_Body_y[1143] = c_Body_y[1142];
                    end else begin
                        n_Body_x[1143] = c_Body_x[c_Size-1];
                        n_Body_y[1143] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1144) begin
                        n_Body_x[1144] = c_Body_x[1143];
                        n_Body_y[1144] = c_Body_y[1143];
                    end else begin
                        n_Body_x[1144] = c_Body_x[c_Size-1];
                        n_Body_y[1144] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1145) begin
                        n_Body_x[1145] = c_Body_x[1144];
                        n_Body_y[1145] = c_Body_y[1144];
                    end else begin
                        n_Body_x[1145] = c_Body_x[c_Size-1];
                        n_Body_y[1145] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1146) begin
                        n_Body_x[1146] = c_Body_x[1145];
                        n_Body_y[1146] = c_Body_y[1145];
                    end else begin
                        n_Body_x[1146] = c_Body_x[c_Size-1];
                        n_Body_y[1146] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1147) begin
                        n_Body_x[1147] = c_Body_x[1146];
                        n_Body_y[1147] = c_Body_y[1146];
                    end else begin
                        n_Body_x[1147] = c_Body_x[c_Size-1];
                        n_Body_y[1147] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1148) begin
                        n_Body_x[1148] = c_Body_x[1147];
                        n_Body_y[1148] = c_Body_y[1147];
                    end else begin
                        n_Body_x[1148] = c_Body_x[c_Size-1];
                        n_Body_y[1148] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1149) begin
                        n_Body_x[1149] = c_Body_x[1148];
                        n_Body_y[1149] = c_Body_y[1148];
                    end else begin
                        n_Body_x[1149] = c_Body_x[c_Size-1];
                        n_Body_y[1149] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1150) begin
                        n_Body_x[1150] = c_Body_x[1149];
                        n_Body_y[1150] = c_Body_y[1149];
                    end else begin
                        n_Body_x[1150] = c_Body_x[c_Size-1];
                        n_Body_y[1150] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1151) begin
                        n_Body_x[1151] = c_Body_x[1150];
                        n_Body_y[1151] = c_Body_y[1150];
                    end else begin
                        n_Body_x[1151] = c_Body_x[c_Size-1];
                        n_Body_y[1151] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1152) begin
                        n_Body_x[1152] = c_Body_x[1151];
                        n_Body_y[1152] = c_Body_y[1151];
                    end else begin
                        n_Body_x[1152] = c_Body_x[c_Size-1];
                        n_Body_y[1152] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1153) begin
                        n_Body_x[1153] = c_Body_x[1152];
                        n_Body_y[1153] = c_Body_y[1152];
                    end else begin
                        n_Body_x[1153] = c_Body_x[c_Size-1];
                        n_Body_y[1153] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1154) begin
                        n_Body_x[1154] = c_Body_x[1153];
                        n_Body_y[1154] = c_Body_y[1153];
                    end else begin
                        n_Body_x[1154] = c_Body_x[c_Size-1];
                        n_Body_y[1154] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1155) begin
                        n_Body_x[1155] = c_Body_x[1154];
                        n_Body_y[1155] = c_Body_y[1154];
                    end else begin
                        n_Body_x[1155] = c_Body_x[c_Size-1];
                        n_Body_y[1155] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1156) begin
                        n_Body_x[1156] = c_Body_x[1155];
                        n_Body_y[1156] = c_Body_y[1155];
                    end else begin
                        n_Body_x[1156] = c_Body_x[c_Size-1];
                        n_Body_y[1156] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1157) begin
                        n_Body_x[1157] = c_Body_x[1156];
                        n_Body_y[1157] = c_Body_y[1156];
                    end else begin
                        n_Body_x[1157] = c_Body_x[c_Size-1];
                        n_Body_y[1157] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1158) begin
                        n_Body_x[1158] = c_Body_x[1157];
                        n_Body_y[1158] = c_Body_y[1157];
                    end else begin
                        n_Body_x[1158] = c_Body_x[c_Size-1];
                        n_Body_y[1158] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1159) begin
                        n_Body_x[1159] = c_Body_x[1158];
                        n_Body_y[1159] = c_Body_y[1158];
                    end else begin
                        n_Body_x[1159] = c_Body_x[c_Size-1];
                        n_Body_y[1159] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1160) begin
                        n_Body_x[1160] = c_Body_x[1159];
                        n_Body_y[1160] = c_Body_y[1159];
                    end else begin
                        n_Body_x[1160] = c_Body_x[c_Size-1];
                        n_Body_y[1160] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1161) begin
                        n_Body_x[1161] = c_Body_x[1160];
                        n_Body_y[1161] = c_Body_y[1160];
                    end else begin
                        n_Body_x[1161] = c_Body_x[c_Size-1];
                        n_Body_y[1161] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1162) begin
                        n_Body_x[1162] = c_Body_x[1161];
                        n_Body_y[1162] = c_Body_y[1161];
                    end else begin
                        n_Body_x[1162] = c_Body_x[c_Size-1];
                        n_Body_y[1162] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1163) begin
                        n_Body_x[1163] = c_Body_x[1162];
                        n_Body_y[1163] = c_Body_y[1162];
                    end else begin
                        n_Body_x[1163] = c_Body_x[c_Size-1];
                        n_Body_y[1163] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1164) begin
                        n_Body_x[1164] = c_Body_x[1163];
                        n_Body_y[1164] = c_Body_y[1163];
                    end else begin
                        n_Body_x[1164] = c_Body_x[c_Size-1];
                        n_Body_y[1164] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1165) begin
                        n_Body_x[1165] = c_Body_x[1164];
                        n_Body_y[1165] = c_Body_y[1164];
                    end else begin
                        n_Body_x[1165] = c_Body_x[c_Size-1];
                        n_Body_y[1165] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1166) begin
                        n_Body_x[1166] = c_Body_x[1165];
                        n_Body_y[1166] = c_Body_y[1165];
                    end else begin
                        n_Body_x[1166] = c_Body_x[c_Size-1];
                        n_Body_y[1166] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1167) begin
                        n_Body_x[1167] = c_Body_x[1166];
                        n_Body_y[1167] = c_Body_y[1166];
                    end else begin
                        n_Body_x[1167] = c_Body_x[c_Size-1];
                        n_Body_y[1167] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1168) begin
                        n_Body_x[1168] = c_Body_x[1167];
                        n_Body_y[1168] = c_Body_y[1167];
                    end else begin
                        n_Body_x[1168] = c_Body_x[c_Size-1];
                        n_Body_y[1168] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1169) begin
                        n_Body_x[1169] = c_Body_x[1168];
                        n_Body_y[1169] = c_Body_y[1168];
                    end else begin
                        n_Body_x[1169] = c_Body_x[c_Size-1];
                        n_Body_y[1169] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1170) begin
                        n_Body_x[1170] = c_Body_x[1169];
                        n_Body_y[1170] = c_Body_y[1169];
                    end else begin
                        n_Body_x[1170] = c_Body_x[c_Size-1];
                        n_Body_y[1170] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1171) begin
                        n_Body_x[1171] = c_Body_x[1170];
                        n_Body_y[1171] = c_Body_y[1170];
                    end else begin
                        n_Body_x[1171] = c_Body_x[c_Size-1];
                        n_Body_y[1171] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1172) begin
                        n_Body_x[1172] = c_Body_x[1171];
                        n_Body_y[1172] = c_Body_y[1171];
                    end else begin
                        n_Body_x[1172] = c_Body_x[c_Size-1];
                        n_Body_y[1172] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1173) begin
                        n_Body_x[1173] = c_Body_x[1172];
                        n_Body_y[1173] = c_Body_y[1172];
                    end else begin
                        n_Body_x[1173] = c_Body_x[c_Size-1];
                        n_Body_y[1173] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1174) begin
                        n_Body_x[1174] = c_Body_x[1173];
                        n_Body_y[1174] = c_Body_y[1173];
                    end else begin
                        n_Body_x[1174] = c_Body_x[c_Size-1];
                        n_Body_y[1174] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1175) begin
                        n_Body_x[1175] = c_Body_x[1174];
                        n_Body_y[1175] = c_Body_y[1174];
                    end else begin
                        n_Body_x[1175] = c_Body_x[c_Size-1];
                        n_Body_y[1175] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1176) begin
                        n_Body_x[1176] = c_Body_x[1175];
                        n_Body_y[1176] = c_Body_y[1175];
                    end else begin
                        n_Body_x[1176] = c_Body_x[c_Size-1];
                        n_Body_y[1176] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1177) begin
                        n_Body_x[1177] = c_Body_x[1176];
                        n_Body_y[1177] = c_Body_y[1176];
                    end else begin
                        n_Body_x[1177] = c_Body_x[c_Size-1];
                        n_Body_y[1177] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1178) begin
                        n_Body_x[1178] = c_Body_x[1177];
                        n_Body_y[1178] = c_Body_y[1177];
                    end else begin
                        n_Body_x[1178] = c_Body_x[c_Size-1];
                        n_Body_y[1178] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1179) begin
                        n_Body_x[1179] = c_Body_x[1178];
                        n_Body_y[1179] = c_Body_y[1178];
                    end else begin
                        n_Body_x[1179] = c_Body_x[c_Size-1];
                        n_Body_y[1179] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1180) begin
                        n_Body_x[1180] = c_Body_x[1179];
                        n_Body_y[1180] = c_Body_y[1179];
                    end else begin
                        n_Body_x[1180] = c_Body_x[c_Size-1];
                        n_Body_y[1180] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1181) begin
                        n_Body_x[1181] = c_Body_x[1180];
                        n_Body_y[1181] = c_Body_y[1180];
                    end else begin
                        n_Body_x[1181] = c_Body_x[c_Size-1];
                        n_Body_y[1181] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1182) begin
                        n_Body_x[1182] = c_Body_x[1181];
                        n_Body_y[1182] = c_Body_y[1181];
                    end else begin
                        n_Body_x[1182] = c_Body_x[c_Size-1];
                        n_Body_y[1182] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1183) begin
                        n_Body_x[1183] = c_Body_x[1182];
                        n_Body_y[1183] = c_Body_y[1182];
                    end else begin
                        n_Body_x[1183] = c_Body_x[c_Size-1];
                        n_Body_y[1183] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1184) begin
                        n_Body_x[1184] = c_Body_x[1183];
                        n_Body_y[1184] = c_Body_y[1183];
                    end else begin
                        n_Body_x[1184] = c_Body_x[c_Size-1];
                        n_Body_y[1184] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1185) begin
                        n_Body_x[1185] = c_Body_x[1184];
                        n_Body_y[1185] = c_Body_y[1184];
                    end else begin
                        n_Body_x[1185] = c_Body_x[c_Size-1];
                        n_Body_y[1185] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1186) begin
                        n_Body_x[1186] = c_Body_x[1185];
                        n_Body_y[1186] = c_Body_y[1185];
                    end else begin
                        n_Body_x[1186] = c_Body_x[c_Size-1];
                        n_Body_y[1186] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1187) begin
                        n_Body_x[1187] = c_Body_x[1186];
                        n_Body_y[1187] = c_Body_y[1186];
                    end else begin
                        n_Body_x[1187] = c_Body_x[c_Size-1];
                        n_Body_y[1187] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1188) begin
                        n_Body_x[1188] = c_Body_x[1187];
                        n_Body_y[1188] = c_Body_y[1187];
                    end else begin
                        n_Body_x[1188] = c_Body_x[c_Size-1];
                        n_Body_y[1188] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1189) begin
                        n_Body_x[1189] = c_Body_x[1188];
                        n_Body_y[1189] = c_Body_y[1188];
                    end else begin
                        n_Body_x[1189] = c_Body_x[c_Size-1];
                        n_Body_y[1189] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1190) begin
                        n_Body_x[1190] = c_Body_x[1189];
                        n_Body_y[1190] = c_Body_y[1189];
                    end else begin
                        n_Body_x[1190] = c_Body_x[c_Size-1];
                        n_Body_y[1190] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1191) begin
                        n_Body_x[1191] = c_Body_x[1190];
                        n_Body_y[1191] = c_Body_y[1190];
                    end else begin
                        n_Body_x[1191] = c_Body_x[c_Size-1];
                        n_Body_y[1191] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1192) begin
                        n_Body_x[1192] = c_Body_x[1191];
                        n_Body_y[1192] = c_Body_y[1191];
                    end else begin
                        n_Body_x[1192] = c_Body_x[c_Size-1];
                        n_Body_y[1192] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1193) begin
                        n_Body_x[1193] = c_Body_x[1192];
                        n_Body_y[1193] = c_Body_y[1192];
                    end else begin
                        n_Body_x[1193] = c_Body_x[c_Size-1];
                        n_Body_y[1193] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1194) begin
                        n_Body_x[1194] = c_Body_x[1193];
                        n_Body_y[1194] = c_Body_y[1193];
                    end else begin
                        n_Body_x[1194] = c_Body_x[c_Size-1];
                        n_Body_y[1194] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1195) begin
                        n_Body_x[1195] = c_Body_x[1194];
                        n_Body_y[1195] = c_Body_y[1194];
                    end else begin
                        n_Body_x[1195] = c_Body_x[c_Size-1];
                        n_Body_y[1195] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1196) begin
                        n_Body_x[1196] = c_Body_x[1195];
                        n_Body_y[1196] = c_Body_y[1195];
                    end else begin
                        n_Body_x[1196] = c_Body_x[c_Size-1];
                        n_Body_y[1196] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1197) begin
                        n_Body_x[1197] = c_Body_x[1196];
                        n_Body_y[1197] = c_Body_y[1196];
                    end else begin
                        n_Body_x[1197] = c_Body_x[c_Size-1];
                        n_Body_y[1197] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1198) begin
                        n_Body_x[1198] = c_Body_x[1197];
                        n_Body_y[1198] = c_Body_y[1197];
                    end else begin
                        n_Body_x[1198] = c_Body_x[c_Size-1];
                        n_Body_y[1198] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1199) begin
                        n_Body_x[1199] = c_Body_x[1198];
                        n_Body_y[1199] = c_Body_y[1198];
                    end else begin
                        n_Body_x[1199] = c_Body_x[c_Size-1];
                        n_Body_y[1199] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1200) begin
                        n_Body_x[1200] = c_Body_x[1199];
                        n_Body_y[1200] = c_Body_y[1199];
                    end else begin
                        n_Body_x[1200] = c_Body_x[c_Size-1];
                        n_Body_y[1200] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1201) begin
                        n_Body_x[1201] = c_Body_x[1200];
                        n_Body_y[1201] = c_Body_y[1200];
                    end else begin
                        n_Body_x[1201] = c_Body_x[c_Size-1];
                        n_Body_y[1201] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1202) begin
                        n_Body_x[1202] = c_Body_x[1201];
                        n_Body_y[1202] = c_Body_y[1201];
                    end else begin
                        n_Body_x[1202] = c_Body_x[c_Size-1];
                        n_Body_y[1202] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1203) begin
                        n_Body_x[1203] = c_Body_x[1202];
                        n_Body_y[1203] = c_Body_y[1202];
                    end else begin
                        n_Body_x[1203] = c_Body_x[c_Size-1];
                        n_Body_y[1203] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1204) begin
                        n_Body_x[1204] = c_Body_x[1203];
                        n_Body_y[1204] = c_Body_y[1203];
                    end else begin
                        n_Body_x[1204] = c_Body_x[c_Size-1];
                        n_Body_y[1204] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1205) begin
                        n_Body_x[1205] = c_Body_x[1204];
                        n_Body_y[1205] = c_Body_y[1204];
                    end else begin
                        n_Body_x[1205] = c_Body_x[c_Size-1];
                        n_Body_y[1205] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1206) begin
                        n_Body_x[1206] = c_Body_x[1205];
                        n_Body_y[1206] = c_Body_y[1205];
                    end else begin
                        n_Body_x[1206] = c_Body_x[c_Size-1];
                        n_Body_y[1206] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1207) begin
                        n_Body_x[1207] = c_Body_x[1206];
                        n_Body_y[1207] = c_Body_y[1206];
                    end else begin
                        n_Body_x[1207] = c_Body_x[c_Size-1];
                        n_Body_y[1207] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1208) begin
                        n_Body_x[1208] = c_Body_x[1207];
                        n_Body_y[1208] = c_Body_y[1207];
                    end else begin
                        n_Body_x[1208] = c_Body_x[c_Size-1];
                        n_Body_y[1208] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1209) begin
                        n_Body_x[1209] = c_Body_x[1208];
                        n_Body_y[1209] = c_Body_y[1208];
                    end else begin
                        n_Body_x[1209] = c_Body_x[c_Size-1];
                        n_Body_y[1209] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1210) begin
                        n_Body_x[1210] = c_Body_x[1209];
                        n_Body_y[1210] = c_Body_y[1209];
                    end else begin
                        n_Body_x[1210] = c_Body_x[c_Size-1];
                        n_Body_y[1210] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1211) begin
                        n_Body_x[1211] = c_Body_x[1210];
                        n_Body_y[1211] = c_Body_y[1210];
                    end else begin
                        n_Body_x[1211] = c_Body_x[c_Size-1];
                        n_Body_y[1211] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1212) begin
                        n_Body_x[1212] = c_Body_x[1211];
                        n_Body_y[1212] = c_Body_y[1211];
                    end else begin
                        n_Body_x[1212] = c_Body_x[c_Size-1];
                        n_Body_y[1212] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1213) begin
                        n_Body_x[1213] = c_Body_x[1212];
                        n_Body_y[1213] = c_Body_y[1212];
                    end else begin
                        n_Body_x[1213] = c_Body_x[c_Size-1];
                        n_Body_y[1213] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1214) begin
                        n_Body_x[1214] = c_Body_x[1213];
                        n_Body_y[1214] = c_Body_y[1213];
                    end else begin
                        n_Body_x[1214] = c_Body_x[c_Size-1];
                        n_Body_y[1214] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1215) begin
                        n_Body_x[1215] = c_Body_x[1214];
                        n_Body_y[1215] = c_Body_y[1214];
                    end else begin
                        n_Body_x[1215] = c_Body_x[c_Size-1];
                        n_Body_y[1215] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1216) begin
                        n_Body_x[1216] = c_Body_x[1215];
                        n_Body_y[1216] = c_Body_y[1215];
                    end else begin
                        n_Body_x[1216] = c_Body_x[c_Size-1];
                        n_Body_y[1216] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1217) begin
                        n_Body_x[1217] = c_Body_x[1216];
                        n_Body_y[1217] = c_Body_y[1216];
                    end else begin
                        n_Body_x[1217] = c_Body_x[c_Size-1];
                        n_Body_y[1217] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1218) begin
                        n_Body_x[1218] = c_Body_x[1217];
                        n_Body_y[1218] = c_Body_y[1217];
                    end else begin
                        n_Body_x[1218] = c_Body_x[c_Size-1];
                        n_Body_y[1218] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1219) begin
                        n_Body_x[1219] = c_Body_x[1218];
                        n_Body_y[1219] = c_Body_y[1218];
                    end else begin
                        n_Body_x[1219] = c_Body_x[c_Size-1];
                        n_Body_y[1219] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1220) begin
                        n_Body_x[1220] = c_Body_x[1219];
                        n_Body_y[1220] = c_Body_y[1219];
                    end else begin
                        n_Body_x[1220] = c_Body_x[c_Size-1];
                        n_Body_y[1220] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1221) begin
                        n_Body_x[1221] = c_Body_x[1220];
                        n_Body_y[1221] = c_Body_y[1220];
                    end else begin
                        n_Body_x[1221] = c_Body_x[c_Size-1];
                        n_Body_y[1221] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1222) begin
                        n_Body_x[1222] = c_Body_x[1221];
                        n_Body_y[1222] = c_Body_y[1221];
                    end else begin
                        n_Body_x[1222] = c_Body_x[c_Size-1];
                        n_Body_y[1222] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1223) begin
                        n_Body_x[1223] = c_Body_x[1222];
                        n_Body_y[1223] = c_Body_y[1222];
                    end else begin
                        n_Body_x[1223] = c_Body_x[c_Size-1];
                        n_Body_y[1223] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1224) begin
                        n_Body_x[1224] = c_Body_x[1223];
                        n_Body_y[1224] = c_Body_y[1223];
                    end else begin
                        n_Body_x[1224] = c_Body_x[c_Size-1];
                        n_Body_y[1224] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1225) begin
                        n_Body_x[1225] = c_Body_x[1224];
                        n_Body_y[1225] = c_Body_y[1224];
                    end else begin
                        n_Body_x[1225] = c_Body_x[c_Size-1];
                        n_Body_y[1225] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1226) begin
                        n_Body_x[1226] = c_Body_x[1225];
                        n_Body_y[1226] = c_Body_y[1225];
                    end else begin
                        n_Body_x[1226] = c_Body_x[c_Size-1];
                        n_Body_y[1226] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1227) begin
                        n_Body_x[1227] = c_Body_x[1226];
                        n_Body_y[1227] = c_Body_y[1226];
                    end else begin
                        n_Body_x[1227] = c_Body_x[c_Size-1];
                        n_Body_y[1227] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1228) begin
                        n_Body_x[1228] = c_Body_x[1227];
                        n_Body_y[1228] = c_Body_y[1227];
                    end else begin
                        n_Body_x[1228] = c_Body_x[c_Size-1];
                        n_Body_y[1228] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1229) begin
                        n_Body_x[1229] = c_Body_x[1228];
                        n_Body_y[1229] = c_Body_y[1228];
                    end else begin
                        n_Body_x[1229] = c_Body_x[c_Size-1];
                        n_Body_y[1229] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1230) begin
                        n_Body_x[1230] = c_Body_x[1229];
                        n_Body_y[1230] = c_Body_y[1229];
                    end else begin
                        n_Body_x[1230] = c_Body_x[c_Size-1];
                        n_Body_y[1230] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1231) begin
                        n_Body_x[1231] = c_Body_x[1230];
                        n_Body_y[1231] = c_Body_y[1230];
                    end else begin
                        n_Body_x[1231] = c_Body_x[c_Size-1];
                        n_Body_y[1231] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1232) begin
                        n_Body_x[1232] = c_Body_x[1231];
                        n_Body_y[1232] = c_Body_y[1231];
                    end else begin
                        n_Body_x[1232] = c_Body_x[c_Size-1];
                        n_Body_y[1232] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1233) begin
                        n_Body_x[1233] = c_Body_x[1232];
                        n_Body_y[1233] = c_Body_y[1232];
                    end else begin
                        n_Body_x[1233] = c_Body_x[c_Size-1];
                        n_Body_y[1233] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1234) begin
                        n_Body_x[1234] = c_Body_x[1233];
                        n_Body_y[1234] = c_Body_y[1233];
                    end else begin
                        n_Body_x[1234] = c_Body_x[c_Size-1];
                        n_Body_y[1234] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1235) begin
                        n_Body_x[1235] = c_Body_x[1234];
                        n_Body_y[1235] = c_Body_y[1234];
                    end else begin
                        n_Body_x[1235] = c_Body_x[c_Size-1];
                        n_Body_y[1235] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1236) begin
                        n_Body_x[1236] = c_Body_x[1235];
                        n_Body_y[1236] = c_Body_y[1235];
                    end else begin
                        n_Body_x[1236] = c_Body_x[c_Size-1];
                        n_Body_y[1236] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1237) begin
                        n_Body_x[1237] = c_Body_x[1236];
                        n_Body_y[1237] = c_Body_y[1236];
                    end else begin
                        n_Body_x[1237] = c_Body_x[c_Size-1];
                        n_Body_y[1237] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1238) begin
                        n_Body_x[1238] = c_Body_x[1237];
                        n_Body_y[1238] = c_Body_y[1237];
                    end else begin
                        n_Body_x[1238] = c_Body_x[c_Size-1];
                        n_Body_y[1238] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1239) begin
                        n_Body_x[1239] = c_Body_x[1238];
                        n_Body_y[1239] = c_Body_y[1238];
                    end else begin
                        n_Body_x[1239] = c_Body_x[c_Size-1];
                        n_Body_y[1239] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1240) begin
                        n_Body_x[1240] = c_Body_x[1239];
                        n_Body_y[1240] = c_Body_y[1239];
                    end else begin
                        n_Body_x[1240] = c_Body_x[c_Size-1];
                        n_Body_y[1240] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1241) begin
                        n_Body_x[1241] = c_Body_x[1240];
                        n_Body_y[1241] = c_Body_y[1240];
                    end else begin
                        n_Body_x[1241] = c_Body_x[c_Size-1];
                        n_Body_y[1241] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1242) begin
                        n_Body_x[1242] = c_Body_x[1241];
                        n_Body_y[1242] = c_Body_y[1241];
                    end else begin
                        n_Body_x[1242] = c_Body_x[c_Size-1];
                        n_Body_y[1242] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1243) begin
                        n_Body_x[1243] = c_Body_x[1242];
                        n_Body_y[1243] = c_Body_y[1242];
                    end else begin
                        n_Body_x[1243] = c_Body_x[c_Size-1];
                        n_Body_y[1243] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1244) begin
                        n_Body_x[1244] = c_Body_x[1243];
                        n_Body_y[1244] = c_Body_y[1243];
                    end else begin
                        n_Body_x[1244] = c_Body_x[c_Size-1];
                        n_Body_y[1244] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1245) begin
                        n_Body_x[1245] = c_Body_x[1244];
                        n_Body_y[1245] = c_Body_y[1244];
                    end else begin
                        n_Body_x[1245] = c_Body_x[c_Size-1];
                        n_Body_y[1245] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1246) begin
                        n_Body_x[1246] = c_Body_x[1245];
                        n_Body_y[1246] = c_Body_y[1245];
                    end else begin
                        n_Body_x[1246] = c_Body_x[c_Size-1];
                        n_Body_y[1246] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1247) begin
                        n_Body_x[1247] = c_Body_x[1246];
                        n_Body_y[1247] = c_Body_y[1246];
                    end else begin
                        n_Body_x[1247] = c_Body_x[c_Size-1];
                        n_Body_y[1247] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1248) begin
                        n_Body_x[1248] = c_Body_x[1247];
                        n_Body_y[1248] = c_Body_y[1247];
                    end else begin
                        n_Body_x[1248] = c_Body_x[c_Size-1];
                        n_Body_y[1248] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1249) begin
                        n_Body_x[1249] = c_Body_x[1248];
                        n_Body_y[1249] = c_Body_y[1248];
                    end else begin
                        n_Body_x[1249] = c_Body_x[c_Size-1];
                        n_Body_y[1249] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1250) begin
                        n_Body_x[1250] = c_Body_x[1249];
                        n_Body_y[1250] = c_Body_y[1249];
                    end else begin
                        n_Body_x[1250] = c_Body_x[c_Size-1];
                        n_Body_y[1250] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1251) begin
                        n_Body_x[1251] = c_Body_x[1250];
                        n_Body_y[1251] = c_Body_y[1250];
                    end else begin
                        n_Body_x[1251] = c_Body_x[c_Size-1];
                        n_Body_y[1251] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1252) begin
                        n_Body_x[1252] = c_Body_x[1251];
                        n_Body_y[1252] = c_Body_y[1251];
                    end else begin
                        n_Body_x[1252] = c_Body_x[c_Size-1];
                        n_Body_y[1252] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1253) begin
                        n_Body_x[1253] = c_Body_x[1252];
                        n_Body_y[1253] = c_Body_y[1252];
                    end else begin
                        n_Body_x[1253] = c_Body_x[c_Size-1];
                        n_Body_y[1253] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1254) begin
                        n_Body_x[1254] = c_Body_x[1253];
                        n_Body_y[1254] = c_Body_y[1253];
                    end else begin
                        n_Body_x[1254] = c_Body_x[c_Size-1];
                        n_Body_y[1254] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1255) begin
                        n_Body_x[1255] = c_Body_x[1254];
                        n_Body_y[1255] = c_Body_y[1254];
                    end else begin
                        n_Body_x[1255] = c_Body_x[c_Size-1];
                        n_Body_y[1255] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1256) begin
                        n_Body_x[1256] = c_Body_x[1255];
                        n_Body_y[1256] = c_Body_y[1255];
                    end else begin
                        n_Body_x[1256] = c_Body_x[c_Size-1];
                        n_Body_y[1256] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1257) begin
                        n_Body_x[1257] = c_Body_x[1256];
                        n_Body_y[1257] = c_Body_y[1256];
                    end else begin
                        n_Body_x[1257] = c_Body_x[c_Size-1];
                        n_Body_y[1257] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1258) begin
                        n_Body_x[1258] = c_Body_x[1257];
                        n_Body_y[1258] = c_Body_y[1257];
                    end else begin
                        n_Body_x[1258] = c_Body_x[c_Size-1];
                        n_Body_y[1258] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1259) begin
                        n_Body_x[1259] = c_Body_x[1258];
                        n_Body_y[1259] = c_Body_y[1258];
                    end else begin
                        n_Body_x[1259] = c_Body_x[c_Size-1];
                        n_Body_y[1259] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1260) begin
                        n_Body_x[1260] = c_Body_x[1259];
                        n_Body_y[1260] = c_Body_y[1259];
                    end else begin
                        n_Body_x[1260] = c_Body_x[c_Size-1];
                        n_Body_y[1260] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1261) begin
                        n_Body_x[1261] = c_Body_x[1260];
                        n_Body_y[1261] = c_Body_y[1260];
                    end else begin
                        n_Body_x[1261] = c_Body_x[c_Size-1];
                        n_Body_y[1261] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1262) begin
                        n_Body_x[1262] = c_Body_x[1261];
                        n_Body_y[1262] = c_Body_y[1261];
                    end else begin
                        n_Body_x[1262] = c_Body_x[c_Size-1];
                        n_Body_y[1262] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1263) begin
                        n_Body_x[1263] = c_Body_x[1262];
                        n_Body_y[1263] = c_Body_y[1262];
                    end else begin
                        n_Body_x[1263] = c_Body_x[c_Size-1];
                        n_Body_y[1263] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1264) begin
                        n_Body_x[1264] = c_Body_x[1263];
                        n_Body_y[1264] = c_Body_y[1263];
                    end else begin
                        n_Body_x[1264] = c_Body_x[c_Size-1];
                        n_Body_y[1264] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1265) begin
                        n_Body_x[1265] = c_Body_x[1264];
                        n_Body_y[1265] = c_Body_y[1264];
                    end else begin
                        n_Body_x[1265] = c_Body_x[c_Size-1];
                        n_Body_y[1265] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1266) begin
                        n_Body_x[1266] = c_Body_x[1265];
                        n_Body_y[1266] = c_Body_y[1265];
                    end else begin
                        n_Body_x[1266] = c_Body_x[c_Size-1];
                        n_Body_y[1266] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1267) begin
                        n_Body_x[1267] = c_Body_x[1266];
                        n_Body_y[1267] = c_Body_y[1266];
                    end else begin
                        n_Body_x[1267] = c_Body_x[c_Size-1];
                        n_Body_y[1267] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1268) begin
                        n_Body_x[1268] = c_Body_x[1267];
                        n_Body_y[1268] = c_Body_y[1267];
                    end else begin
                        n_Body_x[1268] = c_Body_x[c_Size-1];
                        n_Body_y[1268] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1269) begin
                        n_Body_x[1269] = c_Body_x[1268];
                        n_Body_y[1269] = c_Body_y[1268];
                    end else begin
                        n_Body_x[1269] = c_Body_x[c_Size-1];
                        n_Body_y[1269] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1270) begin
                        n_Body_x[1270] = c_Body_x[1269];
                        n_Body_y[1270] = c_Body_y[1269];
                    end else begin
                        n_Body_x[1270] = c_Body_x[c_Size-1];
                        n_Body_y[1270] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1271) begin
                        n_Body_x[1271] = c_Body_x[1270];
                        n_Body_y[1271] = c_Body_y[1270];
                    end else begin
                        n_Body_x[1271] = c_Body_x[c_Size-1];
                        n_Body_y[1271] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1272) begin
                        n_Body_x[1272] = c_Body_x[1271];
                        n_Body_y[1272] = c_Body_y[1271];
                    end else begin
                        n_Body_x[1272] = c_Body_x[c_Size-1];
                        n_Body_y[1272] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1273) begin
                        n_Body_x[1273] = c_Body_x[1272];
                        n_Body_y[1273] = c_Body_y[1272];
                    end else begin
                        n_Body_x[1273] = c_Body_x[c_Size-1];
                        n_Body_y[1273] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1274) begin
                        n_Body_x[1274] = c_Body_x[1273];
                        n_Body_y[1274] = c_Body_y[1273];
                    end else begin
                        n_Body_x[1274] = c_Body_x[c_Size-1];
                        n_Body_y[1274] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1275) begin
                        n_Body_x[1275] = c_Body_x[1274];
                        n_Body_y[1275] = c_Body_y[1274];
                    end else begin
                        n_Body_x[1275] = c_Body_x[c_Size-1];
                        n_Body_y[1275] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1276) begin
                        n_Body_x[1276] = c_Body_x[1275];
                        n_Body_y[1276] = c_Body_y[1275];
                    end else begin
                        n_Body_x[1276] = c_Body_x[c_Size-1];
                        n_Body_y[1276] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1277) begin
                        n_Body_x[1277] = c_Body_x[1276];
                        n_Body_y[1277] = c_Body_y[1276];
                    end else begin
                        n_Body_x[1277] = c_Body_x[c_Size-1];
                        n_Body_y[1277] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1278) begin
                        n_Body_x[1278] = c_Body_x[1277];
                        n_Body_y[1278] = c_Body_y[1277];
                    end else begin
                        n_Body_x[1278] = c_Body_x[c_Size-1];
                        n_Body_y[1278] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1279) begin
                        n_Body_x[1279] = c_Body_x[1278];
                        n_Body_y[1279] = c_Body_y[1278];
                    end else begin
                        n_Body_x[1279] = c_Body_x[c_Size-1];
                        n_Body_y[1279] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1280) begin
                        n_Body_x[1280] = c_Body_x[1279];
                        n_Body_y[1280] = c_Body_y[1279];
                    end else begin
                        n_Body_x[1280] = c_Body_x[c_Size-1];
                        n_Body_y[1280] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1281) begin
                        n_Body_x[1281] = c_Body_x[1280];
                        n_Body_y[1281] = c_Body_y[1280];
                    end else begin
                        n_Body_x[1281] = c_Body_x[c_Size-1];
                        n_Body_y[1281] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1282) begin
                        n_Body_x[1282] = c_Body_x[1281];
                        n_Body_y[1282] = c_Body_y[1281];
                    end else begin
                        n_Body_x[1282] = c_Body_x[c_Size-1];
                        n_Body_y[1282] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1283) begin
                        n_Body_x[1283] = c_Body_x[1282];
                        n_Body_y[1283] = c_Body_y[1282];
                    end else begin
                        n_Body_x[1283] = c_Body_x[c_Size-1];
                        n_Body_y[1283] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1284) begin
                        n_Body_x[1284] = c_Body_x[1283];
                        n_Body_y[1284] = c_Body_y[1283];
                    end else begin
                        n_Body_x[1284] = c_Body_x[c_Size-1];
                        n_Body_y[1284] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1285) begin
                        n_Body_x[1285] = c_Body_x[1284];
                        n_Body_y[1285] = c_Body_y[1284];
                    end else begin
                        n_Body_x[1285] = c_Body_x[c_Size-1];
                        n_Body_y[1285] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1286) begin
                        n_Body_x[1286] = c_Body_x[1285];
                        n_Body_y[1286] = c_Body_y[1285];
                    end else begin
                        n_Body_x[1286] = c_Body_x[c_Size-1];
                        n_Body_y[1286] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1287) begin
                        n_Body_x[1287] = c_Body_x[1286];
                        n_Body_y[1287] = c_Body_y[1286];
                    end else begin
                        n_Body_x[1287] = c_Body_x[c_Size-1];
                        n_Body_y[1287] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1288) begin
                        n_Body_x[1288] = c_Body_x[1287];
                        n_Body_y[1288] = c_Body_y[1287];
                    end else begin
                        n_Body_x[1288] = c_Body_x[c_Size-1];
                        n_Body_y[1288] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1289) begin
                        n_Body_x[1289] = c_Body_x[1288];
                        n_Body_y[1289] = c_Body_y[1288];
                    end else begin
                        n_Body_x[1289] = c_Body_x[c_Size-1];
                        n_Body_y[1289] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1290) begin
                        n_Body_x[1290] = c_Body_x[1289];
                        n_Body_y[1290] = c_Body_y[1289];
                    end else begin
                        n_Body_x[1290] = c_Body_x[c_Size-1];
                        n_Body_y[1290] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1291) begin
                        n_Body_x[1291] = c_Body_x[1290];
                        n_Body_y[1291] = c_Body_y[1290];
                    end else begin
                        n_Body_x[1291] = c_Body_x[c_Size-1];
                        n_Body_y[1291] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1292) begin
                        n_Body_x[1292] = c_Body_x[1291];
                        n_Body_y[1292] = c_Body_y[1291];
                    end else begin
                        n_Body_x[1292] = c_Body_x[c_Size-1];
                        n_Body_y[1292] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1293) begin
                        n_Body_x[1293] = c_Body_x[1292];
                        n_Body_y[1293] = c_Body_y[1292];
                    end else begin
                        n_Body_x[1293] = c_Body_x[c_Size-1];
                        n_Body_y[1293] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1294) begin
                        n_Body_x[1294] = c_Body_x[1293];
                        n_Body_y[1294] = c_Body_y[1293];
                    end else begin
                        n_Body_x[1294] = c_Body_x[c_Size-1];
                        n_Body_y[1294] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1295) begin
                        n_Body_x[1295] = c_Body_x[1294];
                        n_Body_y[1295] = c_Body_y[1294];
                    end else begin
                        n_Body_x[1295] = c_Body_x[c_Size-1];
                        n_Body_y[1295] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1296) begin
                        n_Body_x[1296] = c_Body_x[1295];
                        n_Body_y[1296] = c_Body_y[1295];
                    end else begin
                        n_Body_x[1296] = c_Body_x[c_Size-1];
                        n_Body_y[1296] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1297) begin
                        n_Body_x[1297] = c_Body_x[1296];
                        n_Body_y[1297] = c_Body_y[1296];
                    end else begin
                        n_Body_x[1297] = c_Body_x[c_Size-1];
                        n_Body_y[1297] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1298) begin
                        n_Body_x[1298] = c_Body_x[1297];
                        n_Body_y[1298] = c_Body_y[1297];
                    end else begin
                        n_Body_x[1298] = c_Body_x[c_Size-1];
                        n_Body_y[1298] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1299) begin
                        n_Body_x[1299] = c_Body_x[1298];
                        n_Body_y[1299] = c_Body_y[1298];
                    end else begin
                        n_Body_x[1299] = c_Body_x[c_Size-1];
                        n_Body_y[1299] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1300) begin
                        n_Body_x[1300] = c_Body_x[1299];
                        n_Body_y[1300] = c_Body_y[1299];
                    end else begin
                        n_Body_x[1300] = c_Body_x[c_Size-1];
                        n_Body_y[1300] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1301) begin
                        n_Body_x[1301] = c_Body_x[1300];
                        n_Body_y[1301] = c_Body_y[1300];
                    end else begin
                        n_Body_x[1301] = c_Body_x[c_Size-1];
                        n_Body_y[1301] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1302) begin
                        n_Body_x[1302] = c_Body_x[1301];
                        n_Body_y[1302] = c_Body_y[1301];
                    end else begin
                        n_Body_x[1302] = c_Body_x[c_Size-1];
                        n_Body_y[1302] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1303) begin
                        n_Body_x[1303] = c_Body_x[1302];
                        n_Body_y[1303] = c_Body_y[1302];
                    end else begin
                        n_Body_x[1303] = c_Body_x[c_Size-1];
                        n_Body_y[1303] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1304) begin
                        n_Body_x[1304] = c_Body_x[1303];
                        n_Body_y[1304] = c_Body_y[1303];
                    end else begin
                        n_Body_x[1304] = c_Body_x[c_Size-1];
                        n_Body_y[1304] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1305) begin
                        n_Body_x[1305] = c_Body_x[1304];
                        n_Body_y[1305] = c_Body_y[1304];
                    end else begin
                        n_Body_x[1305] = c_Body_x[c_Size-1];
                        n_Body_y[1305] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1306) begin
                        n_Body_x[1306] = c_Body_x[1305];
                        n_Body_y[1306] = c_Body_y[1305];
                    end else begin
                        n_Body_x[1306] = c_Body_x[c_Size-1];
                        n_Body_y[1306] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1307) begin
                        n_Body_x[1307] = c_Body_x[1306];
                        n_Body_y[1307] = c_Body_y[1306];
                    end else begin
                        n_Body_x[1307] = c_Body_x[c_Size-1];
                        n_Body_y[1307] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1308) begin
                        n_Body_x[1308] = c_Body_x[1307];
                        n_Body_y[1308] = c_Body_y[1307];
                    end else begin
                        n_Body_x[1308] = c_Body_x[c_Size-1];
                        n_Body_y[1308] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1309) begin
                        n_Body_x[1309] = c_Body_x[1308];
                        n_Body_y[1309] = c_Body_y[1308];
                    end else begin
                        n_Body_x[1309] = c_Body_x[c_Size-1];
                        n_Body_y[1309] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1310) begin
                        n_Body_x[1310] = c_Body_x[1309];
                        n_Body_y[1310] = c_Body_y[1309];
                    end else begin
                        n_Body_x[1310] = c_Body_x[c_Size-1];
                        n_Body_y[1310] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1311) begin
                        n_Body_x[1311] = c_Body_x[1310];
                        n_Body_y[1311] = c_Body_y[1310];
                    end else begin
                        n_Body_x[1311] = c_Body_x[c_Size-1];
                        n_Body_y[1311] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1312) begin
                        n_Body_x[1312] = c_Body_x[1311];
                        n_Body_y[1312] = c_Body_y[1311];
                    end else begin
                        n_Body_x[1312] = c_Body_x[c_Size-1];
                        n_Body_y[1312] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1313) begin
                        n_Body_x[1313] = c_Body_x[1312];
                        n_Body_y[1313] = c_Body_y[1312];
                    end else begin
                        n_Body_x[1313] = c_Body_x[c_Size-1];
                        n_Body_y[1313] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1314) begin
                        n_Body_x[1314] = c_Body_x[1313];
                        n_Body_y[1314] = c_Body_y[1313];
                    end else begin
                        n_Body_x[1314] = c_Body_x[c_Size-1];
                        n_Body_y[1314] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1315) begin
                        n_Body_x[1315] = c_Body_x[1314];
                        n_Body_y[1315] = c_Body_y[1314];
                    end else begin
                        n_Body_x[1315] = c_Body_x[c_Size-1];
                        n_Body_y[1315] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1316) begin
                        n_Body_x[1316] = c_Body_x[1315];
                        n_Body_y[1316] = c_Body_y[1315];
                    end else begin
                        n_Body_x[1316] = c_Body_x[c_Size-1];
                        n_Body_y[1316] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1317) begin
                        n_Body_x[1317] = c_Body_x[1316];
                        n_Body_y[1317] = c_Body_y[1316];
                    end else begin
                        n_Body_x[1317] = c_Body_x[c_Size-1];
                        n_Body_y[1317] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1318) begin
                        n_Body_x[1318] = c_Body_x[1317];
                        n_Body_y[1318] = c_Body_y[1317];
                    end else begin
                        n_Body_x[1318] = c_Body_x[c_Size-1];
                        n_Body_y[1318] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1319) begin
                        n_Body_x[1319] = c_Body_x[1318];
                        n_Body_y[1319] = c_Body_y[1318];
                    end else begin
                        n_Body_x[1319] = c_Body_x[c_Size-1];
                        n_Body_y[1319] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1320) begin
                        n_Body_x[1320] = c_Body_x[1319];
                        n_Body_y[1320] = c_Body_y[1319];
                    end else begin
                        n_Body_x[1320] = c_Body_x[c_Size-1];
                        n_Body_y[1320] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1321) begin
                        n_Body_x[1321] = c_Body_x[1320];
                        n_Body_y[1321] = c_Body_y[1320];
                    end else begin
                        n_Body_x[1321] = c_Body_x[c_Size-1];
                        n_Body_y[1321] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1322) begin
                        n_Body_x[1322] = c_Body_x[1321];
                        n_Body_y[1322] = c_Body_y[1321];
                    end else begin
                        n_Body_x[1322] = c_Body_x[c_Size-1];
                        n_Body_y[1322] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1323) begin
                        n_Body_x[1323] = c_Body_x[1322];
                        n_Body_y[1323] = c_Body_y[1322];
                    end else begin
                        n_Body_x[1323] = c_Body_x[c_Size-1];
                        n_Body_y[1323] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1324) begin
                        n_Body_x[1324] = c_Body_x[1323];
                        n_Body_y[1324] = c_Body_y[1323];
                    end else begin
                        n_Body_x[1324] = c_Body_x[c_Size-1];
                        n_Body_y[1324] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1325) begin
                        n_Body_x[1325] = c_Body_x[1324];
                        n_Body_y[1325] = c_Body_y[1324];
                    end else begin
                        n_Body_x[1325] = c_Body_x[c_Size-1];
                        n_Body_y[1325] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1326) begin
                        n_Body_x[1326] = c_Body_x[1325];
                        n_Body_y[1326] = c_Body_y[1325];
                    end else begin
                        n_Body_x[1326] = c_Body_x[c_Size-1];
                        n_Body_y[1326] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1327) begin
                        n_Body_x[1327] = c_Body_x[1326];
                        n_Body_y[1327] = c_Body_y[1326];
                    end else begin
                        n_Body_x[1327] = c_Body_x[c_Size-1];
                        n_Body_y[1327] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1328) begin
                        n_Body_x[1328] = c_Body_x[1327];
                        n_Body_y[1328] = c_Body_y[1327];
                    end else begin
                        n_Body_x[1328] = c_Body_x[c_Size-1];
                        n_Body_y[1328] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1329) begin
                        n_Body_x[1329] = c_Body_x[1328];
                        n_Body_y[1329] = c_Body_y[1328];
                    end else begin
                        n_Body_x[1329] = c_Body_x[c_Size-1];
                        n_Body_y[1329] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1330) begin
                        n_Body_x[1330] = c_Body_x[1329];
                        n_Body_y[1330] = c_Body_y[1329];
                    end else begin
                        n_Body_x[1330] = c_Body_x[c_Size-1];
                        n_Body_y[1330] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1331) begin
                        n_Body_x[1331] = c_Body_x[1330];
                        n_Body_y[1331] = c_Body_y[1330];
                    end else begin
                        n_Body_x[1331] = c_Body_x[c_Size-1];
                        n_Body_y[1331] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1332) begin
                        n_Body_x[1332] = c_Body_x[1331];
                        n_Body_y[1332] = c_Body_y[1331];
                    end else begin
                        n_Body_x[1332] = c_Body_x[c_Size-1];
                        n_Body_y[1332] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1333) begin
                        n_Body_x[1333] = c_Body_x[1332];
                        n_Body_y[1333] = c_Body_y[1332];
                    end else begin
                        n_Body_x[1333] = c_Body_x[c_Size-1];
                        n_Body_y[1333] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1334) begin
                        n_Body_x[1334] = c_Body_x[1333];
                        n_Body_y[1334] = c_Body_y[1333];
                    end else begin
                        n_Body_x[1334] = c_Body_x[c_Size-1];
                        n_Body_y[1334] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1335) begin
                        n_Body_x[1335] = c_Body_x[1334];
                        n_Body_y[1335] = c_Body_y[1334];
                    end else begin
                        n_Body_x[1335] = c_Body_x[c_Size-1];
                        n_Body_y[1335] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1336) begin
                        n_Body_x[1336] = c_Body_x[1335];
                        n_Body_y[1336] = c_Body_y[1335];
                    end else begin
                        n_Body_x[1336] = c_Body_x[c_Size-1];
                        n_Body_y[1336] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1337) begin
                        n_Body_x[1337] = c_Body_x[1336];
                        n_Body_y[1337] = c_Body_y[1336];
                    end else begin
                        n_Body_x[1337] = c_Body_x[c_Size-1];
                        n_Body_y[1337] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1338) begin
                        n_Body_x[1338] = c_Body_x[1337];
                        n_Body_y[1338] = c_Body_y[1337];
                    end else begin
                        n_Body_x[1338] = c_Body_x[c_Size-1];
                        n_Body_y[1338] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1339) begin
                        n_Body_x[1339] = c_Body_x[1338];
                        n_Body_y[1339] = c_Body_y[1338];
                    end else begin
                        n_Body_x[1339] = c_Body_x[c_Size-1];
                        n_Body_y[1339] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1340) begin
                        n_Body_x[1340] = c_Body_x[1339];
                        n_Body_y[1340] = c_Body_y[1339];
                    end else begin
                        n_Body_x[1340] = c_Body_x[c_Size-1];
                        n_Body_y[1340] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1341) begin
                        n_Body_x[1341] = c_Body_x[1340];
                        n_Body_y[1341] = c_Body_y[1340];
                    end else begin
                        n_Body_x[1341] = c_Body_x[c_Size-1];
                        n_Body_y[1341] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1342) begin
                        n_Body_x[1342] = c_Body_x[1341];
                        n_Body_y[1342] = c_Body_y[1341];
                    end else begin
                        n_Body_x[1342] = c_Body_x[c_Size-1];
                        n_Body_y[1342] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1343) begin
                        n_Body_x[1343] = c_Body_x[1342];
                        n_Body_y[1343] = c_Body_y[1342];
                    end else begin
                        n_Body_x[1343] = c_Body_x[c_Size-1];
                        n_Body_y[1343] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1344) begin
                        n_Body_x[1344] = c_Body_x[1343];
                        n_Body_y[1344] = c_Body_y[1343];
                    end else begin
                        n_Body_x[1344] = c_Body_x[c_Size-1];
                        n_Body_y[1344] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1345) begin
                        n_Body_x[1345] = c_Body_x[1344];
                        n_Body_y[1345] = c_Body_y[1344];
                    end else begin
                        n_Body_x[1345] = c_Body_x[c_Size-1];
                        n_Body_y[1345] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1346) begin
                        n_Body_x[1346] = c_Body_x[1345];
                        n_Body_y[1346] = c_Body_y[1345];
                    end else begin
                        n_Body_x[1346] = c_Body_x[c_Size-1];
                        n_Body_y[1346] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1347) begin
                        n_Body_x[1347] = c_Body_x[1346];
                        n_Body_y[1347] = c_Body_y[1346];
                    end else begin
                        n_Body_x[1347] = c_Body_x[c_Size-1];
                        n_Body_y[1347] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1348) begin
                        n_Body_x[1348] = c_Body_x[1347];
                        n_Body_y[1348] = c_Body_y[1347];
                    end else begin
                        n_Body_x[1348] = c_Body_x[c_Size-1];
                        n_Body_y[1348] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1349) begin
                        n_Body_x[1349] = c_Body_x[1348];
                        n_Body_y[1349] = c_Body_y[1348];
                    end else begin
                        n_Body_x[1349] = c_Body_x[c_Size-1];
                        n_Body_y[1349] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1350) begin
                        n_Body_x[1350] = c_Body_x[1349];
                        n_Body_y[1350] = c_Body_y[1349];
                    end else begin
                        n_Body_x[1350] = c_Body_x[c_Size-1];
                        n_Body_y[1350] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1351) begin
                        n_Body_x[1351] = c_Body_x[1350];
                        n_Body_y[1351] = c_Body_y[1350];
                    end else begin
                        n_Body_x[1351] = c_Body_x[c_Size-1];
                        n_Body_y[1351] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1352) begin
                        n_Body_x[1352] = c_Body_x[1351];
                        n_Body_y[1352] = c_Body_y[1351];
                    end else begin
                        n_Body_x[1352] = c_Body_x[c_Size-1];
                        n_Body_y[1352] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1353) begin
                        n_Body_x[1353] = c_Body_x[1352];
                        n_Body_y[1353] = c_Body_y[1352];
                    end else begin
                        n_Body_x[1353] = c_Body_x[c_Size-1];
                        n_Body_y[1353] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1354) begin
                        n_Body_x[1354] = c_Body_x[1353];
                        n_Body_y[1354] = c_Body_y[1353];
                    end else begin
                        n_Body_x[1354] = c_Body_x[c_Size-1];
                        n_Body_y[1354] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1355) begin
                        n_Body_x[1355] = c_Body_x[1354];
                        n_Body_y[1355] = c_Body_y[1354];
                    end else begin
                        n_Body_x[1355] = c_Body_x[c_Size-1];
                        n_Body_y[1355] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1356) begin
                        n_Body_x[1356] = c_Body_x[1355];
                        n_Body_y[1356] = c_Body_y[1355];
                    end else begin
                        n_Body_x[1356] = c_Body_x[c_Size-1];
                        n_Body_y[1356] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1357) begin
                        n_Body_x[1357] = c_Body_x[1356];
                        n_Body_y[1357] = c_Body_y[1356];
                    end else begin
                        n_Body_x[1357] = c_Body_x[c_Size-1];
                        n_Body_y[1357] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1358) begin
                        n_Body_x[1358] = c_Body_x[1357];
                        n_Body_y[1358] = c_Body_y[1357];
                    end else begin
                        n_Body_x[1358] = c_Body_x[c_Size-1];
                        n_Body_y[1358] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1359) begin
                        n_Body_x[1359] = c_Body_x[1358];
                        n_Body_y[1359] = c_Body_y[1358];
                    end else begin
                        n_Body_x[1359] = c_Body_x[c_Size-1];
                        n_Body_y[1359] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1360) begin
                        n_Body_x[1360] = c_Body_x[1359];
                        n_Body_y[1360] = c_Body_y[1359];
                    end else begin
                        n_Body_x[1360] = c_Body_x[c_Size-1];
                        n_Body_y[1360] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1361) begin
                        n_Body_x[1361] = c_Body_x[1360];
                        n_Body_y[1361] = c_Body_y[1360];
                    end else begin
                        n_Body_x[1361] = c_Body_x[c_Size-1];
                        n_Body_y[1361] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1362) begin
                        n_Body_x[1362] = c_Body_x[1361];
                        n_Body_y[1362] = c_Body_y[1361];
                    end else begin
                        n_Body_x[1362] = c_Body_x[c_Size-1];
                        n_Body_y[1362] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1363) begin
                        n_Body_x[1363] = c_Body_x[1362];
                        n_Body_y[1363] = c_Body_y[1362];
                    end else begin
                        n_Body_x[1363] = c_Body_x[c_Size-1];
                        n_Body_y[1363] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1364) begin
                        n_Body_x[1364] = c_Body_x[1363];
                        n_Body_y[1364] = c_Body_y[1363];
                    end else begin
                        n_Body_x[1364] = c_Body_x[c_Size-1];
                        n_Body_y[1364] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1365) begin
                        n_Body_x[1365] = c_Body_x[1364];
                        n_Body_y[1365] = c_Body_y[1364];
                    end else begin
                        n_Body_x[1365] = c_Body_x[c_Size-1];
                        n_Body_y[1365] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1366) begin
                        n_Body_x[1366] = c_Body_x[1365];
                        n_Body_y[1366] = c_Body_y[1365];
                    end else begin
                        n_Body_x[1366] = c_Body_x[c_Size-1];
                        n_Body_y[1366] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1367) begin
                        n_Body_x[1367] = c_Body_x[1366];
                        n_Body_y[1367] = c_Body_y[1366];
                    end else begin
                        n_Body_x[1367] = c_Body_x[c_Size-1];
                        n_Body_y[1367] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1368) begin
                        n_Body_x[1368] = c_Body_x[1367];
                        n_Body_y[1368] = c_Body_y[1367];
                    end else begin
                        n_Body_x[1368] = c_Body_x[c_Size-1];
                        n_Body_y[1368] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1369) begin
                        n_Body_x[1369] = c_Body_x[1368];
                        n_Body_y[1369] = c_Body_y[1368];
                    end else begin
                        n_Body_x[1369] = c_Body_x[c_Size-1];
                        n_Body_y[1369] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1370) begin
                        n_Body_x[1370] = c_Body_x[1369];
                        n_Body_y[1370] = c_Body_y[1369];
                    end else begin
                        n_Body_x[1370] = c_Body_x[c_Size-1];
                        n_Body_y[1370] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1371) begin
                        n_Body_x[1371] = c_Body_x[1370];
                        n_Body_y[1371] = c_Body_y[1370];
                    end else begin
                        n_Body_x[1371] = c_Body_x[c_Size-1];
                        n_Body_y[1371] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1372) begin
                        n_Body_x[1372] = c_Body_x[1371];
                        n_Body_y[1372] = c_Body_y[1371];
                    end else begin
                        n_Body_x[1372] = c_Body_x[c_Size-1];
                        n_Body_y[1372] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1373) begin
                        n_Body_x[1373] = c_Body_x[1372];
                        n_Body_y[1373] = c_Body_y[1372];
                    end else begin
                        n_Body_x[1373] = c_Body_x[c_Size-1];
                        n_Body_y[1373] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1374) begin
                        n_Body_x[1374] = c_Body_x[1373];
                        n_Body_y[1374] = c_Body_y[1373];
                    end else begin
                        n_Body_x[1374] = c_Body_x[c_Size-1];
                        n_Body_y[1374] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1375) begin
                        n_Body_x[1375] = c_Body_x[1374];
                        n_Body_y[1375] = c_Body_y[1374];
                    end else begin
                        n_Body_x[1375] = c_Body_x[c_Size-1];
                        n_Body_y[1375] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1376) begin
                        n_Body_x[1376] = c_Body_x[1375];
                        n_Body_y[1376] = c_Body_y[1375];
                    end else begin
                        n_Body_x[1376] = c_Body_x[c_Size-1];
                        n_Body_y[1376] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1377) begin
                        n_Body_x[1377] = c_Body_x[1376];
                        n_Body_y[1377] = c_Body_y[1376];
                    end else begin
                        n_Body_x[1377] = c_Body_x[c_Size-1];
                        n_Body_y[1377] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1378) begin
                        n_Body_x[1378] = c_Body_x[1377];
                        n_Body_y[1378] = c_Body_y[1377];
                    end else begin
                        n_Body_x[1378] = c_Body_x[c_Size-1];
                        n_Body_y[1378] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1379) begin
                        n_Body_x[1379] = c_Body_x[1378];
                        n_Body_y[1379] = c_Body_y[1378];
                    end else begin
                        n_Body_x[1379] = c_Body_x[c_Size-1];
                        n_Body_y[1379] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1380) begin
                        n_Body_x[1380] = c_Body_x[1379];
                        n_Body_y[1380] = c_Body_y[1379];
                    end else begin
                        n_Body_x[1380] = c_Body_x[c_Size-1];
                        n_Body_y[1380] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1381) begin
                        n_Body_x[1381] = c_Body_x[1380];
                        n_Body_y[1381] = c_Body_y[1380];
                    end else begin
                        n_Body_x[1381] = c_Body_x[c_Size-1];
                        n_Body_y[1381] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1382) begin
                        n_Body_x[1382] = c_Body_x[1381];
                        n_Body_y[1382] = c_Body_y[1381];
                    end else begin
                        n_Body_x[1382] = c_Body_x[c_Size-1];
                        n_Body_y[1382] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1383) begin
                        n_Body_x[1383] = c_Body_x[1382];
                        n_Body_y[1383] = c_Body_y[1382];
                    end else begin
                        n_Body_x[1383] = c_Body_x[c_Size-1];
                        n_Body_y[1383] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1384) begin
                        n_Body_x[1384] = c_Body_x[1383];
                        n_Body_y[1384] = c_Body_y[1383];
                    end else begin
                        n_Body_x[1384] = c_Body_x[c_Size-1];
                        n_Body_y[1384] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1385) begin
                        n_Body_x[1385] = c_Body_x[1384];
                        n_Body_y[1385] = c_Body_y[1384];
                    end else begin
                        n_Body_x[1385] = c_Body_x[c_Size-1];
                        n_Body_y[1385] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1386) begin
                        n_Body_x[1386] = c_Body_x[1385];
                        n_Body_y[1386] = c_Body_y[1385];
                    end else begin
                        n_Body_x[1386] = c_Body_x[c_Size-1];
                        n_Body_y[1386] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1387) begin
                        n_Body_x[1387] = c_Body_x[1386];
                        n_Body_y[1387] = c_Body_y[1386];
                    end else begin
                        n_Body_x[1387] = c_Body_x[c_Size-1];
                        n_Body_y[1387] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1388) begin
                        n_Body_x[1388] = c_Body_x[1387];
                        n_Body_y[1388] = c_Body_y[1387];
                    end else begin
                        n_Body_x[1388] = c_Body_x[c_Size-1];
                        n_Body_y[1388] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1389) begin
                        n_Body_x[1389] = c_Body_x[1388];
                        n_Body_y[1389] = c_Body_y[1388];
                    end else begin
                        n_Body_x[1389] = c_Body_x[c_Size-1];
                        n_Body_y[1389] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1390) begin
                        n_Body_x[1390] = c_Body_x[1389];
                        n_Body_y[1390] = c_Body_y[1389];
                    end else begin
                        n_Body_x[1390] = c_Body_x[c_Size-1];
                        n_Body_y[1390] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1391) begin
                        n_Body_x[1391] = c_Body_x[1390];
                        n_Body_y[1391] = c_Body_y[1390];
                    end else begin
                        n_Body_x[1391] = c_Body_x[c_Size-1];
                        n_Body_y[1391] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1392) begin
                        n_Body_x[1392] = c_Body_x[1391];
                        n_Body_y[1392] = c_Body_y[1391];
                    end else begin
                        n_Body_x[1392] = c_Body_x[c_Size-1];
                        n_Body_y[1392] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1393) begin
                        n_Body_x[1393] = c_Body_x[1392];
                        n_Body_y[1393] = c_Body_y[1392];
                    end else begin
                        n_Body_x[1393] = c_Body_x[c_Size-1];
                        n_Body_y[1393] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1394) begin
                        n_Body_x[1394] = c_Body_x[1393];
                        n_Body_y[1394] = c_Body_y[1393];
                    end else begin
                        n_Body_x[1394] = c_Body_x[c_Size-1];
                        n_Body_y[1394] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1395) begin
                        n_Body_x[1395] = c_Body_x[1394];
                        n_Body_y[1395] = c_Body_y[1394];
                    end else begin
                        n_Body_x[1395] = c_Body_x[c_Size-1];
                        n_Body_y[1395] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1396) begin
                        n_Body_x[1396] = c_Body_x[1395];
                        n_Body_y[1396] = c_Body_y[1395];
                    end else begin
                        n_Body_x[1396] = c_Body_x[c_Size-1];
                        n_Body_y[1396] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1397) begin
                        n_Body_x[1397] = c_Body_x[1396];
                        n_Body_y[1397] = c_Body_y[1396];
                    end else begin
                        n_Body_x[1397] = c_Body_x[c_Size-1];
                        n_Body_y[1397] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1398) begin
                        n_Body_x[1398] = c_Body_x[1397];
                        n_Body_y[1398] = c_Body_y[1397];
                    end else begin
                        n_Body_x[1398] = c_Body_x[c_Size-1];
                        n_Body_y[1398] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1399) begin
                        n_Body_x[1399] = c_Body_x[1398];
                        n_Body_y[1399] = c_Body_y[1398];
                    end else begin
                        n_Body_x[1399] = c_Body_x[c_Size-1];
                        n_Body_y[1399] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1400) begin
                        n_Body_x[1400] = c_Body_x[1399];
                        n_Body_y[1400] = c_Body_y[1399];
                    end else begin
                        n_Body_x[1400] = c_Body_x[c_Size-1];
                        n_Body_y[1400] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1401) begin
                        n_Body_x[1401] = c_Body_x[1400];
                        n_Body_y[1401] = c_Body_y[1400];
                    end else begin
                        n_Body_x[1401] = c_Body_x[c_Size-1];
                        n_Body_y[1401] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1402) begin
                        n_Body_x[1402] = c_Body_x[1401];
                        n_Body_y[1402] = c_Body_y[1401];
                    end else begin
                        n_Body_x[1402] = c_Body_x[c_Size-1];
                        n_Body_y[1402] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1403) begin
                        n_Body_x[1403] = c_Body_x[1402];
                        n_Body_y[1403] = c_Body_y[1402];
                    end else begin
                        n_Body_x[1403] = c_Body_x[c_Size-1];
                        n_Body_y[1403] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1404) begin
                        n_Body_x[1404] = c_Body_x[1403];
                        n_Body_y[1404] = c_Body_y[1403];
                    end else begin
                        n_Body_x[1404] = c_Body_x[c_Size-1];
                        n_Body_y[1404] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1405) begin
                        n_Body_x[1405] = c_Body_x[1404];
                        n_Body_y[1405] = c_Body_y[1404];
                    end else begin
                        n_Body_x[1405] = c_Body_x[c_Size-1];
                        n_Body_y[1405] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1406) begin
                        n_Body_x[1406] = c_Body_x[1405];
                        n_Body_y[1406] = c_Body_y[1405];
                    end else begin
                        n_Body_x[1406] = c_Body_x[c_Size-1];
                        n_Body_y[1406] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1407) begin
                        n_Body_x[1407] = c_Body_x[1406];
                        n_Body_y[1407] = c_Body_y[1406];
                    end else begin
                        n_Body_x[1407] = c_Body_x[c_Size-1];
                        n_Body_y[1407] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1408) begin
                        n_Body_x[1408] = c_Body_x[1407];
                        n_Body_y[1408] = c_Body_y[1407];
                    end else begin
                        n_Body_x[1408] = c_Body_x[c_Size-1];
                        n_Body_y[1408] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1409) begin
                        n_Body_x[1409] = c_Body_x[1408];
                        n_Body_y[1409] = c_Body_y[1408];
                    end else begin
                        n_Body_x[1409] = c_Body_x[c_Size-1];
                        n_Body_y[1409] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1410) begin
                        n_Body_x[1410] = c_Body_x[1409];
                        n_Body_y[1410] = c_Body_y[1409];
                    end else begin
                        n_Body_x[1410] = c_Body_x[c_Size-1];
                        n_Body_y[1410] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1411) begin
                        n_Body_x[1411] = c_Body_x[1410];
                        n_Body_y[1411] = c_Body_y[1410];
                    end else begin
                        n_Body_x[1411] = c_Body_x[c_Size-1];
                        n_Body_y[1411] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1412) begin
                        n_Body_x[1412] = c_Body_x[1411];
                        n_Body_y[1412] = c_Body_y[1411];
                    end else begin
                        n_Body_x[1412] = c_Body_x[c_Size-1];
                        n_Body_y[1412] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1413) begin
                        n_Body_x[1413] = c_Body_x[1412];
                        n_Body_y[1413] = c_Body_y[1412];
                    end else begin
                        n_Body_x[1413] = c_Body_x[c_Size-1];
                        n_Body_y[1413] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1414) begin
                        n_Body_x[1414] = c_Body_x[1413];
                        n_Body_y[1414] = c_Body_y[1413];
                    end else begin
                        n_Body_x[1414] = c_Body_x[c_Size-1];
                        n_Body_y[1414] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1415) begin
                        n_Body_x[1415] = c_Body_x[1414];
                        n_Body_y[1415] = c_Body_y[1414];
                    end else begin
                        n_Body_x[1415] = c_Body_x[c_Size-1];
                        n_Body_y[1415] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1416) begin
                        n_Body_x[1416] = c_Body_x[1415];
                        n_Body_y[1416] = c_Body_y[1415];
                    end else begin
                        n_Body_x[1416] = c_Body_x[c_Size-1];
                        n_Body_y[1416] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1417) begin
                        n_Body_x[1417] = c_Body_x[1416];
                        n_Body_y[1417] = c_Body_y[1416];
                    end else begin
                        n_Body_x[1417] = c_Body_x[c_Size-1];
                        n_Body_y[1417] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1418) begin
                        n_Body_x[1418] = c_Body_x[1417];
                        n_Body_y[1418] = c_Body_y[1417];
                    end else begin
                        n_Body_x[1418] = c_Body_x[c_Size-1];
                        n_Body_y[1418] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1419) begin
                        n_Body_x[1419] = c_Body_x[1418];
                        n_Body_y[1419] = c_Body_y[1418];
                    end else begin
                        n_Body_x[1419] = c_Body_x[c_Size-1];
                        n_Body_y[1419] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1420) begin
                        n_Body_x[1420] = c_Body_x[1419];
                        n_Body_y[1420] = c_Body_y[1419];
                    end else begin
                        n_Body_x[1420] = c_Body_x[c_Size-1];
                        n_Body_y[1420] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1421) begin
                        n_Body_x[1421] = c_Body_x[1420];
                        n_Body_y[1421] = c_Body_y[1420];
                    end else begin
                        n_Body_x[1421] = c_Body_x[c_Size-1];
                        n_Body_y[1421] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1422) begin
                        n_Body_x[1422] = c_Body_x[1421];
                        n_Body_y[1422] = c_Body_y[1421];
                    end else begin
                        n_Body_x[1422] = c_Body_x[c_Size-1];
                        n_Body_y[1422] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1423) begin
                        n_Body_x[1423] = c_Body_x[1422];
                        n_Body_y[1423] = c_Body_y[1422];
                    end else begin
                        n_Body_x[1423] = c_Body_x[c_Size-1];
                        n_Body_y[1423] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1424) begin
                        n_Body_x[1424] = c_Body_x[1423];
                        n_Body_y[1424] = c_Body_y[1423];
                    end else begin
                        n_Body_x[1424] = c_Body_x[c_Size-1];
                        n_Body_y[1424] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1425) begin
                        n_Body_x[1425] = c_Body_x[1424];
                        n_Body_y[1425] = c_Body_y[1424];
                    end else begin
                        n_Body_x[1425] = c_Body_x[c_Size-1];
                        n_Body_y[1425] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1426) begin
                        n_Body_x[1426] = c_Body_x[1425];
                        n_Body_y[1426] = c_Body_y[1425];
                    end else begin
                        n_Body_x[1426] = c_Body_x[c_Size-1];
                        n_Body_y[1426] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1427) begin
                        n_Body_x[1427] = c_Body_x[1426];
                        n_Body_y[1427] = c_Body_y[1426];
                    end else begin
                        n_Body_x[1427] = c_Body_x[c_Size-1];
                        n_Body_y[1427] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1428) begin
                        n_Body_x[1428] = c_Body_x[1427];
                        n_Body_y[1428] = c_Body_y[1427];
                    end else begin
                        n_Body_x[1428] = c_Body_x[c_Size-1];
                        n_Body_y[1428] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1429) begin
                        n_Body_x[1429] = c_Body_x[1428];
                        n_Body_y[1429] = c_Body_y[1428];
                    end else begin
                        n_Body_x[1429] = c_Body_x[c_Size-1];
                        n_Body_y[1429] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1430) begin
                        n_Body_x[1430] = c_Body_x[1429];
                        n_Body_y[1430] = c_Body_y[1429];
                    end else begin
                        n_Body_x[1430] = c_Body_x[c_Size-1];
                        n_Body_y[1430] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1431) begin
                        n_Body_x[1431] = c_Body_x[1430];
                        n_Body_y[1431] = c_Body_y[1430];
                    end else begin
                        n_Body_x[1431] = c_Body_x[c_Size-1];
                        n_Body_y[1431] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1432) begin
                        n_Body_x[1432] = c_Body_x[1431];
                        n_Body_y[1432] = c_Body_y[1431];
                    end else begin
                        n_Body_x[1432] = c_Body_x[c_Size-1];
                        n_Body_y[1432] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1433) begin
                        n_Body_x[1433] = c_Body_x[1432];
                        n_Body_y[1433] = c_Body_y[1432];
                    end else begin
                        n_Body_x[1433] = c_Body_x[c_Size-1];
                        n_Body_y[1433] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1434) begin
                        n_Body_x[1434] = c_Body_x[1433];
                        n_Body_y[1434] = c_Body_y[1433];
                    end else begin
                        n_Body_x[1434] = c_Body_x[c_Size-1];
                        n_Body_y[1434] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1435) begin
                        n_Body_x[1435] = c_Body_x[1434];
                        n_Body_y[1435] = c_Body_y[1434];
                    end else begin
                        n_Body_x[1435] = c_Body_x[c_Size-1];
                        n_Body_y[1435] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1436) begin
                        n_Body_x[1436] = c_Body_x[1435];
                        n_Body_y[1436] = c_Body_y[1435];
                    end else begin
                        n_Body_x[1436] = c_Body_x[c_Size-1];
                        n_Body_y[1436] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1437) begin
                        n_Body_x[1437] = c_Body_x[1436];
                        n_Body_y[1437] = c_Body_y[1436];
                    end else begin
                        n_Body_x[1437] = c_Body_x[c_Size-1];
                        n_Body_y[1437] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1438) begin
                        n_Body_x[1438] = c_Body_x[1437];
                        n_Body_y[1438] = c_Body_y[1437];
                    end else begin
                        n_Body_x[1438] = c_Body_x[c_Size-1];
                        n_Body_y[1438] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1439) begin
                        n_Body_x[1439] = c_Body_x[1438];
                        n_Body_y[1439] = c_Body_y[1438];
                    end else begin
                        n_Body_x[1439] = c_Body_x[c_Size-1];
                        n_Body_y[1439] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1440) begin
                        n_Body_x[1440] = c_Body_x[1439];
                        n_Body_y[1440] = c_Body_y[1439];
                    end else begin
                        n_Body_x[1440] = c_Body_x[c_Size-1];
                        n_Body_y[1440] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1441) begin
                        n_Body_x[1441] = c_Body_x[1440];
                        n_Body_y[1441] = c_Body_y[1440];
                    end else begin
                        n_Body_x[1441] = c_Body_x[c_Size-1];
                        n_Body_y[1441] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1442) begin
                        n_Body_x[1442] = c_Body_x[1441];
                        n_Body_y[1442] = c_Body_y[1441];
                    end else begin
                        n_Body_x[1442] = c_Body_x[c_Size-1];
                        n_Body_y[1442] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1443) begin
                        n_Body_x[1443] = c_Body_x[1442];
                        n_Body_y[1443] = c_Body_y[1442];
                    end else begin
                        n_Body_x[1443] = c_Body_x[c_Size-1];
                        n_Body_y[1443] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1444) begin
                        n_Body_x[1444] = c_Body_x[1443];
                        n_Body_y[1444] = c_Body_y[1443];
                    end else begin
                        n_Body_x[1444] = c_Body_x[c_Size-1];
                        n_Body_y[1444] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1445) begin
                        n_Body_x[1445] = c_Body_x[1444];
                        n_Body_y[1445] = c_Body_y[1444];
                    end else begin
                        n_Body_x[1445] = c_Body_x[c_Size-1];
                        n_Body_y[1445] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1446) begin
                        n_Body_x[1446] = c_Body_x[1445];
                        n_Body_y[1446] = c_Body_y[1445];
                    end else begin
                        n_Body_x[1446] = c_Body_x[c_Size-1];
                        n_Body_y[1446] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1447) begin
                        n_Body_x[1447] = c_Body_x[1446];
                        n_Body_y[1447] = c_Body_y[1446];
                    end else begin
                        n_Body_x[1447] = c_Body_x[c_Size-1];
                        n_Body_y[1447] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1448) begin
                        n_Body_x[1448] = c_Body_x[1447];
                        n_Body_y[1448] = c_Body_y[1447];
                    end else begin
                        n_Body_x[1448] = c_Body_x[c_Size-1];
                        n_Body_y[1448] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1449) begin
                        n_Body_x[1449] = c_Body_x[1448];
                        n_Body_y[1449] = c_Body_y[1448];
                    end else begin
                        n_Body_x[1449] = c_Body_x[c_Size-1];
                        n_Body_y[1449] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1450) begin
                        n_Body_x[1450] = c_Body_x[1449];
                        n_Body_y[1450] = c_Body_y[1449];
                    end else begin
                        n_Body_x[1450] = c_Body_x[c_Size-1];
                        n_Body_y[1450] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1451) begin
                        n_Body_x[1451] = c_Body_x[1450];
                        n_Body_y[1451] = c_Body_y[1450];
                    end else begin
                        n_Body_x[1451] = c_Body_x[c_Size-1];
                        n_Body_y[1451] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1452) begin
                        n_Body_x[1452] = c_Body_x[1451];
                        n_Body_y[1452] = c_Body_y[1451];
                    end else begin
                        n_Body_x[1452] = c_Body_x[c_Size-1];
                        n_Body_y[1452] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1453) begin
                        n_Body_x[1453] = c_Body_x[1452];
                        n_Body_y[1453] = c_Body_y[1452];
                    end else begin
                        n_Body_x[1453] = c_Body_x[c_Size-1];
                        n_Body_y[1453] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1454) begin
                        n_Body_x[1454] = c_Body_x[1453];
                        n_Body_y[1454] = c_Body_y[1453];
                    end else begin
                        n_Body_x[1454] = c_Body_x[c_Size-1];
                        n_Body_y[1454] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1455) begin
                        n_Body_x[1455] = c_Body_x[1454];
                        n_Body_y[1455] = c_Body_y[1454];
                    end else begin
                        n_Body_x[1455] = c_Body_x[c_Size-1];
                        n_Body_y[1455] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1456) begin
                        n_Body_x[1456] = c_Body_x[1455];
                        n_Body_y[1456] = c_Body_y[1455];
                    end else begin
                        n_Body_x[1456] = c_Body_x[c_Size-1];
                        n_Body_y[1456] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1457) begin
                        n_Body_x[1457] = c_Body_x[1456];
                        n_Body_y[1457] = c_Body_y[1456];
                    end else begin
                        n_Body_x[1457] = c_Body_x[c_Size-1];
                        n_Body_y[1457] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1458) begin
                        n_Body_x[1458] = c_Body_x[1457];
                        n_Body_y[1458] = c_Body_y[1457];
                    end else begin
                        n_Body_x[1458] = c_Body_x[c_Size-1];
                        n_Body_y[1458] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1459) begin
                        n_Body_x[1459] = c_Body_x[1458];
                        n_Body_y[1459] = c_Body_y[1458];
                    end else begin
                        n_Body_x[1459] = c_Body_x[c_Size-1];
                        n_Body_y[1459] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1460) begin
                        n_Body_x[1460] = c_Body_x[1459];
                        n_Body_y[1460] = c_Body_y[1459];
                    end else begin
                        n_Body_x[1460] = c_Body_x[c_Size-1];
                        n_Body_y[1460] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1461) begin
                        n_Body_x[1461] = c_Body_x[1460];
                        n_Body_y[1461] = c_Body_y[1460];
                    end else begin
                        n_Body_x[1461] = c_Body_x[c_Size-1];
                        n_Body_y[1461] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1462) begin
                        n_Body_x[1462] = c_Body_x[1461];
                        n_Body_y[1462] = c_Body_y[1461];
                    end else begin
                        n_Body_x[1462] = c_Body_x[c_Size-1];
                        n_Body_y[1462] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1463) begin
                        n_Body_x[1463] = c_Body_x[1462];
                        n_Body_y[1463] = c_Body_y[1462];
                    end else begin
                        n_Body_x[1463] = c_Body_x[c_Size-1];
                        n_Body_y[1463] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1464) begin
                        n_Body_x[1464] = c_Body_x[1463];
                        n_Body_y[1464] = c_Body_y[1463];
                    end else begin
                        n_Body_x[1464] = c_Body_x[c_Size-1];
                        n_Body_y[1464] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1465) begin
                        n_Body_x[1465] = c_Body_x[1464];
                        n_Body_y[1465] = c_Body_y[1464];
                    end else begin
                        n_Body_x[1465] = c_Body_x[c_Size-1];
                        n_Body_y[1465] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1466) begin
                        n_Body_x[1466] = c_Body_x[1465];
                        n_Body_y[1466] = c_Body_y[1465];
                    end else begin
                        n_Body_x[1466] = c_Body_x[c_Size-1];
                        n_Body_y[1466] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1467) begin
                        n_Body_x[1467] = c_Body_x[1466];
                        n_Body_y[1467] = c_Body_y[1466];
                    end else begin
                        n_Body_x[1467] = c_Body_x[c_Size-1];
                        n_Body_y[1467] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1468) begin
                        n_Body_x[1468] = c_Body_x[1467];
                        n_Body_y[1468] = c_Body_y[1467];
                    end else begin
                        n_Body_x[1468] = c_Body_x[c_Size-1];
                        n_Body_y[1468] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1469) begin
                        n_Body_x[1469] = c_Body_x[1468];
                        n_Body_y[1469] = c_Body_y[1468];
                    end else begin
                        n_Body_x[1469] = c_Body_x[c_Size-1];
                        n_Body_y[1469] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1470) begin
                        n_Body_x[1470] = c_Body_x[1469];
                        n_Body_y[1470] = c_Body_y[1469];
                    end else begin
                        n_Body_x[1470] = c_Body_x[c_Size-1];
                        n_Body_y[1470] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1471) begin
                        n_Body_x[1471] = c_Body_x[1470];
                        n_Body_y[1471] = c_Body_y[1470];
                    end else begin
                        n_Body_x[1471] = c_Body_x[c_Size-1];
                        n_Body_y[1471] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1472) begin
                        n_Body_x[1472] = c_Body_x[1471];
                        n_Body_y[1472] = c_Body_y[1471];
                    end else begin
                        n_Body_x[1472] = c_Body_x[c_Size-1];
                        n_Body_y[1472] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1473) begin
                        n_Body_x[1473] = c_Body_x[1472];
                        n_Body_y[1473] = c_Body_y[1472];
                    end else begin
                        n_Body_x[1473] = c_Body_x[c_Size-1];
                        n_Body_y[1473] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1474) begin
                        n_Body_x[1474] = c_Body_x[1473];
                        n_Body_y[1474] = c_Body_y[1473];
                    end else begin
                        n_Body_x[1474] = c_Body_x[c_Size-1];
                        n_Body_y[1474] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1475) begin
                        n_Body_x[1475] = c_Body_x[1474];
                        n_Body_y[1475] = c_Body_y[1474];
                    end else begin
                        n_Body_x[1475] = c_Body_x[c_Size-1];
                        n_Body_y[1475] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1476) begin
                        n_Body_x[1476] = c_Body_x[1475];
                        n_Body_y[1476] = c_Body_y[1475];
                    end else begin
                        n_Body_x[1476] = c_Body_x[c_Size-1];
                        n_Body_y[1476] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1477) begin
                        n_Body_x[1477] = c_Body_x[1476];
                        n_Body_y[1477] = c_Body_y[1476];
                    end else begin
                        n_Body_x[1477] = c_Body_x[c_Size-1];
                        n_Body_y[1477] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1478) begin
                        n_Body_x[1478] = c_Body_x[1477];
                        n_Body_y[1478] = c_Body_y[1477];
                    end else begin
                        n_Body_x[1478] = c_Body_x[c_Size-1];
                        n_Body_y[1478] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1479) begin
                        n_Body_x[1479] = c_Body_x[1478];
                        n_Body_y[1479] = c_Body_y[1478];
                    end else begin
                        n_Body_x[1479] = c_Body_x[c_Size-1];
                        n_Body_y[1479] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1480) begin
                        n_Body_x[1480] = c_Body_x[1479];
                        n_Body_y[1480] = c_Body_y[1479];
                    end else begin
                        n_Body_x[1480] = c_Body_x[c_Size-1];
                        n_Body_y[1480] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1481) begin
                        n_Body_x[1481] = c_Body_x[1480];
                        n_Body_y[1481] = c_Body_y[1480];
                    end else begin
                        n_Body_x[1481] = c_Body_x[c_Size-1];
                        n_Body_y[1481] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1482) begin
                        n_Body_x[1482] = c_Body_x[1481];
                        n_Body_y[1482] = c_Body_y[1481];
                    end else begin
                        n_Body_x[1482] = c_Body_x[c_Size-1];
                        n_Body_y[1482] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1483) begin
                        n_Body_x[1483] = c_Body_x[1482];
                        n_Body_y[1483] = c_Body_y[1482];
                    end else begin
                        n_Body_x[1483] = c_Body_x[c_Size-1];
                        n_Body_y[1483] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1484) begin
                        n_Body_x[1484] = c_Body_x[1483];
                        n_Body_y[1484] = c_Body_y[1483];
                    end else begin
                        n_Body_x[1484] = c_Body_x[c_Size-1];
                        n_Body_y[1484] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1485) begin
                        n_Body_x[1485] = c_Body_x[1484];
                        n_Body_y[1485] = c_Body_y[1484];
                    end else begin
                        n_Body_x[1485] = c_Body_x[c_Size-1];
                        n_Body_y[1485] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1486) begin
                        n_Body_x[1486] = c_Body_x[1485];
                        n_Body_y[1486] = c_Body_y[1485];
                    end else begin
                        n_Body_x[1486] = c_Body_x[c_Size-1];
                        n_Body_y[1486] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1487) begin
                        n_Body_x[1487] = c_Body_x[1486];
                        n_Body_y[1487] = c_Body_y[1486];
                    end else begin
                        n_Body_x[1487] = c_Body_x[c_Size-1];
                        n_Body_y[1487] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1488) begin
                        n_Body_x[1488] = c_Body_x[1487];
                        n_Body_y[1488] = c_Body_y[1487];
                    end else begin
                        n_Body_x[1488] = c_Body_x[c_Size-1];
                        n_Body_y[1488] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1489) begin
                        n_Body_x[1489] = c_Body_x[1488];
                        n_Body_y[1489] = c_Body_y[1488];
                    end else begin
                        n_Body_x[1489] = c_Body_x[c_Size-1];
                        n_Body_y[1489] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1490) begin
                        n_Body_x[1490] = c_Body_x[1489];
                        n_Body_y[1490] = c_Body_y[1489];
                    end else begin
                        n_Body_x[1490] = c_Body_x[c_Size-1];
                        n_Body_y[1490] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1491) begin
                        n_Body_x[1491] = c_Body_x[1490];
                        n_Body_y[1491] = c_Body_y[1490];
                    end else begin
                        n_Body_x[1491] = c_Body_x[c_Size-1];
                        n_Body_y[1491] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1492) begin
                        n_Body_x[1492] = c_Body_x[1491];
                        n_Body_y[1492] = c_Body_y[1491];
                    end else begin
                        n_Body_x[1492] = c_Body_x[c_Size-1];
                        n_Body_y[1492] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1493) begin
                        n_Body_x[1493] = c_Body_x[1492];
                        n_Body_y[1493] = c_Body_y[1492];
                    end else begin
                        n_Body_x[1493] = c_Body_x[c_Size-1];
                        n_Body_y[1493] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1494) begin
                        n_Body_x[1494] = c_Body_x[1493];
                        n_Body_y[1494] = c_Body_y[1493];
                    end else begin
                        n_Body_x[1494] = c_Body_x[c_Size-1];
                        n_Body_y[1494] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1495) begin
                        n_Body_x[1495] = c_Body_x[1494];
                        n_Body_y[1495] = c_Body_y[1494];
                    end else begin
                        n_Body_x[1495] = c_Body_x[c_Size-1];
                        n_Body_y[1495] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1496) begin
                        n_Body_x[1496] = c_Body_x[1495];
                        n_Body_y[1496] = c_Body_y[1495];
                    end else begin
                        n_Body_x[1496] = c_Body_x[c_Size-1];
                        n_Body_y[1496] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1497) begin
                        n_Body_x[1497] = c_Body_x[1496];
                        n_Body_y[1497] = c_Body_y[1496];
                    end else begin
                        n_Body_x[1497] = c_Body_x[c_Size-1];
                        n_Body_y[1497] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1498) begin
                        n_Body_x[1498] = c_Body_x[1497];
                        n_Body_y[1498] = c_Body_y[1497];
                    end else begin
                        n_Body_x[1498] = c_Body_x[c_Size-1];
                        n_Body_y[1498] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1499) begin
                        n_Body_x[1499] = c_Body_x[1498];
                        n_Body_y[1499] = c_Body_y[1498];
                    end else begin
                        n_Body_x[1499] = c_Body_x[c_Size-1];
                        n_Body_y[1499] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1500) begin
                        n_Body_x[1500] = c_Body_x[1499];
                        n_Body_y[1500] = c_Body_y[1499];
                    end else begin
                        n_Body_x[1500] = c_Body_x[c_Size-1];
                        n_Body_y[1500] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1501) begin
                        n_Body_x[1501] = c_Body_x[1500];
                        n_Body_y[1501] = c_Body_y[1500];
                    end else begin
                        n_Body_x[1501] = c_Body_x[c_Size-1];
                        n_Body_y[1501] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1502) begin
                        n_Body_x[1502] = c_Body_x[1501];
                        n_Body_y[1502] = c_Body_y[1501];
                    end else begin
                        n_Body_x[1502] = c_Body_x[c_Size-1];
                        n_Body_y[1502] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1503) begin
                        n_Body_x[1503] = c_Body_x[1502];
                        n_Body_y[1503] = c_Body_y[1502];
                    end else begin
                        n_Body_x[1503] = c_Body_x[c_Size-1];
                        n_Body_y[1503] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1504) begin
                        n_Body_x[1504] = c_Body_x[1503];
                        n_Body_y[1504] = c_Body_y[1503];
                    end else begin
                        n_Body_x[1504] = c_Body_x[c_Size-1];
                        n_Body_y[1504] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1505) begin
                        n_Body_x[1505] = c_Body_x[1504];
                        n_Body_y[1505] = c_Body_y[1504];
                    end else begin
                        n_Body_x[1505] = c_Body_x[c_Size-1];
                        n_Body_y[1505] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1506) begin
                        n_Body_x[1506] = c_Body_x[1505];
                        n_Body_y[1506] = c_Body_y[1505];
                    end else begin
                        n_Body_x[1506] = c_Body_x[c_Size-1];
                        n_Body_y[1506] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1507) begin
                        n_Body_x[1507] = c_Body_x[1506];
                        n_Body_y[1507] = c_Body_y[1506];
                    end else begin
                        n_Body_x[1507] = c_Body_x[c_Size-1];
                        n_Body_y[1507] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1508) begin
                        n_Body_x[1508] = c_Body_x[1507];
                        n_Body_y[1508] = c_Body_y[1507];
                    end else begin
                        n_Body_x[1508] = c_Body_x[c_Size-1];
                        n_Body_y[1508] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1509) begin
                        n_Body_x[1509] = c_Body_x[1508];
                        n_Body_y[1509] = c_Body_y[1508];
                    end else begin
                        n_Body_x[1509] = c_Body_x[c_Size-1];
                        n_Body_y[1509] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1510) begin
                        n_Body_x[1510] = c_Body_x[1509];
                        n_Body_y[1510] = c_Body_y[1509];
                    end else begin
                        n_Body_x[1510] = c_Body_x[c_Size-1];
                        n_Body_y[1510] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1511) begin
                        n_Body_x[1511] = c_Body_x[1510];
                        n_Body_y[1511] = c_Body_y[1510];
                    end else begin
                        n_Body_x[1511] = c_Body_x[c_Size-1];
                        n_Body_y[1511] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1512) begin
                        n_Body_x[1512] = c_Body_x[1511];
                        n_Body_y[1512] = c_Body_y[1511];
                    end else begin
                        n_Body_x[1512] = c_Body_x[c_Size-1];
                        n_Body_y[1512] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1513) begin
                        n_Body_x[1513] = c_Body_x[1512];
                        n_Body_y[1513] = c_Body_y[1512];
                    end else begin
                        n_Body_x[1513] = c_Body_x[c_Size-1];
                        n_Body_y[1513] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1514) begin
                        n_Body_x[1514] = c_Body_x[1513];
                        n_Body_y[1514] = c_Body_y[1513];
                    end else begin
                        n_Body_x[1514] = c_Body_x[c_Size-1];
                        n_Body_y[1514] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1515) begin
                        n_Body_x[1515] = c_Body_x[1514];
                        n_Body_y[1515] = c_Body_y[1514];
                    end else begin
                        n_Body_x[1515] = c_Body_x[c_Size-1];
                        n_Body_y[1515] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1516) begin
                        n_Body_x[1516] = c_Body_x[1515];
                        n_Body_y[1516] = c_Body_y[1515];
                    end else begin
                        n_Body_x[1516] = c_Body_x[c_Size-1];
                        n_Body_y[1516] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1517) begin
                        n_Body_x[1517] = c_Body_x[1516];
                        n_Body_y[1517] = c_Body_y[1516];
                    end else begin
                        n_Body_x[1517] = c_Body_x[c_Size-1];
                        n_Body_y[1517] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1518) begin
                        n_Body_x[1518] = c_Body_x[1517];
                        n_Body_y[1518] = c_Body_y[1517];
                    end else begin
                        n_Body_x[1518] = c_Body_x[c_Size-1];
                        n_Body_y[1518] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1519) begin
                        n_Body_x[1519] = c_Body_x[1518];
                        n_Body_y[1519] = c_Body_y[1518];
                    end else begin
                        n_Body_x[1519] = c_Body_x[c_Size-1];
                        n_Body_y[1519] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1520) begin
                        n_Body_x[1520] = c_Body_x[1519];
                        n_Body_y[1520] = c_Body_y[1519];
                    end else begin
                        n_Body_x[1520] = c_Body_x[c_Size-1];
                        n_Body_y[1520] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1521) begin
                        n_Body_x[1521] = c_Body_x[1520];
                        n_Body_y[1521] = c_Body_y[1520];
                    end else begin
                        n_Body_x[1521] = c_Body_x[c_Size-1];
                        n_Body_y[1521] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1522) begin
                        n_Body_x[1522] = c_Body_x[1521];
                        n_Body_y[1522] = c_Body_y[1521];
                    end else begin
                        n_Body_x[1522] = c_Body_x[c_Size-1];
                        n_Body_y[1522] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1523) begin
                        n_Body_x[1523] = c_Body_x[1522];
                        n_Body_y[1523] = c_Body_y[1522];
                    end else begin
                        n_Body_x[1523] = c_Body_x[c_Size-1];
                        n_Body_y[1523] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1524) begin
                        n_Body_x[1524] = c_Body_x[1523];
                        n_Body_y[1524] = c_Body_y[1523];
                    end else begin
                        n_Body_x[1524] = c_Body_x[c_Size-1];
                        n_Body_y[1524] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1525) begin
                        n_Body_x[1525] = c_Body_x[1524];
                        n_Body_y[1525] = c_Body_y[1524];
                    end else begin
                        n_Body_x[1525] = c_Body_x[c_Size-1];
                        n_Body_y[1525] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1526) begin
                        n_Body_x[1526] = c_Body_x[1525];
                        n_Body_y[1526] = c_Body_y[1525];
                    end else begin
                        n_Body_x[1526] = c_Body_x[c_Size-1];
                        n_Body_y[1526] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1527) begin
                        n_Body_x[1527] = c_Body_x[1526];
                        n_Body_y[1527] = c_Body_y[1526];
                    end else begin
                        n_Body_x[1527] = c_Body_x[c_Size-1];
                        n_Body_y[1527] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1528) begin
                        n_Body_x[1528] = c_Body_x[1527];
                        n_Body_y[1528] = c_Body_y[1527];
                    end else begin
                        n_Body_x[1528] = c_Body_x[c_Size-1];
                        n_Body_y[1528] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1529) begin
                        n_Body_x[1529] = c_Body_x[1528];
                        n_Body_y[1529] = c_Body_y[1528];
                    end else begin
                        n_Body_x[1529] = c_Body_x[c_Size-1];
                        n_Body_y[1529] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1530) begin
                        n_Body_x[1530] = c_Body_x[1529];
                        n_Body_y[1530] = c_Body_y[1529];
                    end else begin
                        n_Body_x[1530] = c_Body_x[c_Size-1];
                        n_Body_y[1530] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1531) begin
                        n_Body_x[1531] = c_Body_x[1530];
                        n_Body_y[1531] = c_Body_y[1530];
                    end else begin
                        n_Body_x[1531] = c_Body_x[c_Size-1];
                        n_Body_y[1531] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1532) begin
                        n_Body_x[1532] = c_Body_x[1531];
                        n_Body_y[1532] = c_Body_y[1531];
                    end else begin
                        n_Body_x[1532] = c_Body_x[c_Size-1];
                        n_Body_y[1532] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1533) begin
                        n_Body_x[1533] = c_Body_x[1532];
                        n_Body_y[1533] = c_Body_y[1532];
                    end else begin
                        n_Body_x[1533] = c_Body_x[c_Size-1];
                        n_Body_y[1533] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1534) begin
                        n_Body_x[1534] = c_Body_x[1533];
                        n_Body_y[1534] = c_Body_y[1533];
                    end else begin
                        n_Body_x[1534] = c_Body_x[c_Size-1];
                        n_Body_y[1534] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1535) begin
                        n_Body_x[1535] = c_Body_x[1534];
                        n_Body_y[1535] = c_Body_y[1534];
                    end else begin
                        n_Body_x[1535] = c_Body_x[c_Size-1];
                        n_Body_y[1535] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1536) begin
                        n_Body_x[1536] = c_Body_x[1535];
                        n_Body_y[1536] = c_Body_y[1535];
                    end else begin
                        n_Body_x[1536] = c_Body_x[c_Size-1];
                        n_Body_y[1536] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1537) begin
                        n_Body_x[1537] = c_Body_x[1536];
                        n_Body_y[1537] = c_Body_y[1536];
                    end else begin
                        n_Body_x[1537] = c_Body_x[c_Size-1];
                        n_Body_y[1537] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1538) begin
                        n_Body_x[1538] = c_Body_x[1537];
                        n_Body_y[1538] = c_Body_y[1537];
                    end else begin
                        n_Body_x[1538] = c_Body_x[c_Size-1];
                        n_Body_y[1538] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1539) begin
                        n_Body_x[1539] = c_Body_x[1538];
                        n_Body_y[1539] = c_Body_y[1538];
                    end else begin
                        n_Body_x[1539] = c_Body_x[c_Size-1];
                        n_Body_y[1539] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1540) begin
                        n_Body_x[1540] = c_Body_x[1539];
                        n_Body_y[1540] = c_Body_y[1539];
                    end else begin
                        n_Body_x[1540] = c_Body_x[c_Size-1];
                        n_Body_y[1540] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1541) begin
                        n_Body_x[1541] = c_Body_x[1540];
                        n_Body_y[1541] = c_Body_y[1540];
                    end else begin
                        n_Body_x[1541] = c_Body_x[c_Size-1];
                        n_Body_y[1541] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1542) begin
                        n_Body_x[1542] = c_Body_x[1541];
                        n_Body_y[1542] = c_Body_y[1541];
                    end else begin
                        n_Body_x[1542] = c_Body_x[c_Size-1];
                        n_Body_y[1542] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1543) begin
                        n_Body_x[1543] = c_Body_x[1542];
                        n_Body_y[1543] = c_Body_y[1542];
                    end else begin
                        n_Body_x[1543] = c_Body_x[c_Size-1];
                        n_Body_y[1543] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1544) begin
                        n_Body_x[1544] = c_Body_x[1543];
                        n_Body_y[1544] = c_Body_y[1543];
                    end else begin
                        n_Body_x[1544] = c_Body_x[c_Size-1];
                        n_Body_y[1544] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1545) begin
                        n_Body_x[1545] = c_Body_x[1544];
                        n_Body_y[1545] = c_Body_y[1544];
                    end else begin
                        n_Body_x[1545] = c_Body_x[c_Size-1];
                        n_Body_y[1545] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1546) begin
                        n_Body_x[1546] = c_Body_x[1545];
                        n_Body_y[1546] = c_Body_y[1545];
                    end else begin
                        n_Body_x[1546] = c_Body_x[c_Size-1];
                        n_Body_y[1546] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1547) begin
                        n_Body_x[1547] = c_Body_x[1546];
                        n_Body_y[1547] = c_Body_y[1546];
                    end else begin
                        n_Body_x[1547] = c_Body_x[c_Size-1];
                        n_Body_y[1547] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1548) begin
                        n_Body_x[1548] = c_Body_x[1547];
                        n_Body_y[1548] = c_Body_y[1547];
                    end else begin
                        n_Body_x[1548] = c_Body_x[c_Size-1];
                        n_Body_y[1548] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1549) begin
                        n_Body_x[1549] = c_Body_x[1548];
                        n_Body_y[1549] = c_Body_y[1548];
                    end else begin
                        n_Body_x[1549] = c_Body_x[c_Size-1];
                        n_Body_y[1549] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1550) begin
                        n_Body_x[1550] = c_Body_x[1549];
                        n_Body_y[1550] = c_Body_y[1549];
                    end else begin
                        n_Body_x[1550] = c_Body_x[c_Size-1];
                        n_Body_y[1550] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1551) begin
                        n_Body_x[1551] = c_Body_x[1550];
                        n_Body_y[1551] = c_Body_y[1550];
                    end else begin
                        n_Body_x[1551] = c_Body_x[c_Size-1];
                        n_Body_y[1551] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1552) begin
                        n_Body_x[1552] = c_Body_x[1551];
                        n_Body_y[1552] = c_Body_y[1551];
                    end else begin
                        n_Body_x[1552] = c_Body_x[c_Size-1];
                        n_Body_y[1552] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1553) begin
                        n_Body_x[1553] = c_Body_x[1552];
                        n_Body_y[1553] = c_Body_y[1552];
                    end else begin
                        n_Body_x[1553] = c_Body_x[c_Size-1];
                        n_Body_y[1553] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1554) begin
                        n_Body_x[1554] = c_Body_x[1553];
                        n_Body_y[1554] = c_Body_y[1553];
                    end else begin
                        n_Body_x[1554] = c_Body_x[c_Size-1];
                        n_Body_y[1554] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1555) begin
                        n_Body_x[1555] = c_Body_x[1554];
                        n_Body_y[1555] = c_Body_y[1554];
                    end else begin
                        n_Body_x[1555] = c_Body_x[c_Size-1];
                        n_Body_y[1555] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1556) begin
                        n_Body_x[1556] = c_Body_x[1555];
                        n_Body_y[1556] = c_Body_y[1555];
                    end else begin
                        n_Body_x[1556] = c_Body_x[c_Size-1];
                        n_Body_y[1556] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1557) begin
                        n_Body_x[1557] = c_Body_x[1556];
                        n_Body_y[1557] = c_Body_y[1556];
                    end else begin
                        n_Body_x[1557] = c_Body_x[c_Size-1];
                        n_Body_y[1557] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1558) begin
                        n_Body_x[1558] = c_Body_x[1557];
                        n_Body_y[1558] = c_Body_y[1557];
                    end else begin
                        n_Body_x[1558] = c_Body_x[c_Size-1];
                        n_Body_y[1558] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1559) begin
                        n_Body_x[1559] = c_Body_x[1558];
                        n_Body_y[1559] = c_Body_y[1558];
                    end else begin
                        n_Body_x[1559] = c_Body_x[c_Size-1];
                        n_Body_y[1559] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1560) begin
                        n_Body_x[1560] = c_Body_x[1559];
                        n_Body_y[1560] = c_Body_y[1559];
                    end else begin
                        n_Body_x[1560] = c_Body_x[c_Size-1];
                        n_Body_y[1560] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1561) begin
                        n_Body_x[1561] = c_Body_x[1560];
                        n_Body_y[1561] = c_Body_y[1560];
                    end else begin
                        n_Body_x[1561] = c_Body_x[c_Size-1];
                        n_Body_y[1561] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1562) begin
                        n_Body_x[1562] = c_Body_x[1561];
                        n_Body_y[1562] = c_Body_y[1561];
                    end else begin
                        n_Body_x[1562] = c_Body_x[c_Size-1];
                        n_Body_y[1562] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1563) begin
                        n_Body_x[1563] = c_Body_x[1562];
                        n_Body_y[1563] = c_Body_y[1562];
                    end else begin
                        n_Body_x[1563] = c_Body_x[c_Size-1];
                        n_Body_y[1563] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1564) begin
                        n_Body_x[1564] = c_Body_x[1563];
                        n_Body_y[1564] = c_Body_y[1563];
                    end else begin
                        n_Body_x[1564] = c_Body_x[c_Size-1];
                        n_Body_y[1564] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1565) begin
                        n_Body_x[1565] = c_Body_x[1564];
                        n_Body_y[1565] = c_Body_y[1564];
                    end else begin
                        n_Body_x[1565] = c_Body_x[c_Size-1];
                        n_Body_y[1565] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1566) begin
                        n_Body_x[1566] = c_Body_x[1565];
                        n_Body_y[1566] = c_Body_y[1565];
                    end else begin
                        n_Body_x[1566] = c_Body_x[c_Size-1];
                        n_Body_y[1566] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1567) begin
                        n_Body_x[1567] = c_Body_x[1566];
                        n_Body_y[1567] = c_Body_y[1566];
                    end else begin
                        n_Body_x[1567] = c_Body_x[c_Size-1];
                        n_Body_y[1567] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1568) begin
                        n_Body_x[1568] = c_Body_x[1567];
                        n_Body_y[1568] = c_Body_y[1567];
                    end else begin
                        n_Body_x[1568] = c_Body_x[c_Size-1];
                        n_Body_y[1568] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1569) begin
                        n_Body_x[1569] = c_Body_x[1568];
                        n_Body_y[1569] = c_Body_y[1568];
                    end else begin
                        n_Body_x[1569] = c_Body_x[c_Size-1];
                        n_Body_y[1569] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1570) begin
                        n_Body_x[1570] = c_Body_x[1569];
                        n_Body_y[1570] = c_Body_y[1569];
                    end else begin
                        n_Body_x[1570] = c_Body_x[c_Size-1];
                        n_Body_y[1570] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1571) begin
                        n_Body_x[1571] = c_Body_x[1570];
                        n_Body_y[1571] = c_Body_y[1570];
                    end else begin
                        n_Body_x[1571] = c_Body_x[c_Size-1];
                        n_Body_y[1571] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1572) begin
                        n_Body_x[1572] = c_Body_x[1571];
                        n_Body_y[1572] = c_Body_y[1571];
                    end else begin
                        n_Body_x[1572] = c_Body_x[c_Size-1];
                        n_Body_y[1572] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1573) begin
                        n_Body_x[1573] = c_Body_x[1572];
                        n_Body_y[1573] = c_Body_y[1572];
                    end else begin
                        n_Body_x[1573] = c_Body_x[c_Size-1];
                        n_Body_y[1573] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1574) begin
                        n_Body_x[1574] = c_Body_x[1573];
                        n_Body_y[1574] = c_Body_y[1573];
                    end else begin
                        n_Body_x[1574] = c_Body_x[c_Size-1];
                        n_Body_y[1574] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1575) begin
                        n_Body_x[1575] = c_Body_x[1574];
                        n_Body_y[1575] = c_Body_y[1574];
                    end else begin
                        n_Body_x[1575] = c_Body_x[c_Size-1];
                        n_Body_y[1575] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1576) begin
                        n_Body_x[1576] = c_Body_x[1575];
                        n_Body_y[1576] = c_Body_y[1575];
                    end else begin
                        n_Body_x[1576] = c_Body_x[c_Size-1];
                        n_Body_y[1576] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1577) begin
                        n_Body_x[1577] = c_Body_x[1576];
                        n_Body_y[1577] = c_Body_y[1576];
                    end else begin
                        n_Body_x[1577] = c_Body_x[c_Size-1];
                        n_Body_y[1577] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1578) begin
                        n_Body_x[1578] = c_Body_x[1577];
                        n_Body_y[1578] = c_Body_y[1577];
                    end else begin
                        n_Body_x[1578] = c_Body_x[c_Size-1];
                        n_Body_y[1578] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1579) begin
                        n_Body_x[1579] = c_Body_x[1578];
                        n_Body_y[1579] = c_Body_y[1578];
                    end else begin
                        n_Body_x[1579] = c_Body_x[c_Size-1];
                        n_Body_y[1579] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1580) begin
                        n_Body_x[1580] = c_Body_x[1579];
                        n_Body_y[1580] = c_Body_y[1579];
                    end else begin
                        n_Body_x[1580] = c_Body_x[c_Size-1];
                        n_Body_y[1580] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1581) begin
                        n_Body_x[1581] = c_Body_x[1580];
                        n_Body_y[1581] = c_Body_y[1580];
                    end else begin
                        n_Body_x[1581] = c_Body_x[c_Size-1];
                        n_Body_y[1581] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1582) begin
                        n_Body_x[1582] = c_Body_x[1581];
                        n_Body_y[1582] = c_Body_y[1581];
                    end else begin
                        n_Body_x[1582] = c_Body_x[c_Size-1];
                        n_Body_y[1582] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1583) begin
                        n_Body_x[1583] = c_Body_x[1582];
                        n_Body_y[1583] = c_Body_y[1582];
                    end else begin
                        n_Body_x[1583] = c_Body_x[c_Size-1];
                        n_Body_y[1583] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1584) begin
                        n_Body_x[1584] = c_Body_x[1583];
                        n_Body_y[1584] = c_Body_y[1583];
                    end else begin
                        n_Body_x[1584] = c_Body_x[c_Size-1];
                        n_Body_y[1584] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1585) begin
                        n_Body_x[1585] = c_Body_x[1584];
                        n_Body_y[1585] = c_Body_y[1584];
                    end else begin
                        n_Body_x[1585] = c_Body_x[c_Size-1];
                        n_Body_y[1585] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1586) begin
                        n_Body_x[1586] = c_Body_x[1585];
                        n_Body_y[1586] = c_Body_y[1585];
                    end else begin
                        n_Body_x[1586] = c_Body_x[c_Size-1];
                        n_Body_y[1586] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1587) begin
                        n_Body_x[1587] = c_Body_x[1586];
                        n_Body_y[1587] = c_Body_y[1586];
                    end else begin
                        n_Body_x[1587] = c_Body_x[c_Size-1];
                        n_Body_y[1587] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1588) begin
                        n_Body_x[1588] = c_Body_x[1587];
                        n_Body_y[1588] = c_Body_y[1587];
                    end else begin
                        n_Body_x[1588] = c_Body_x[c_Size-1];
                        n_Body_y[1588] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1589) begin
                        n_Body_x[1589] = c_Body_x[1588];
                        n_Body_y[1589] = c_Body_y[1588];
                    end else begin
                        n_Body_x[1589] = c_Body_x[c_Size-1];
                        n_Body_y[1589] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1590) begin
                        n_Body_x[1590] = c_Body_x[1589];
                        n_Body_y[1590] = c_Body_y[1589];
                    end else begin
                        n_Body_x[1590] = c_Body_x[c_Size-1];
                        n_Body_y[1590] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1591) begin
                        n_Body_x[1591] = c_Body_x[1590];
                        n_Body_y[1591] = c_Body_y[1590];
                    end else begin
                        n_Body_x[1591] = c_Body_x[c_Size-1];
                        n_Body_y[1591] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1592) begin
                        n_Body_x[1592] = c_Body_x[1591];
                        n_Body_y[1592] = c_Body_y[1591];
                    end else begin
                        n_Body_x[1592] = c_Body_x[c_Size-1];
                        n_Body_y[1592] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1593) begin
                        n_Body_x[1593] = c_Body_x[1592];
                        n_Body_y[1593] = c_Body_y[1592];
                    end else begin
                        n_Body_x[1593] = c_Body_x[c_Size-1];
                        n_Body_y[1593] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1594) begin
                        n_Body_x[1594] = c_Body_x[1593];
                        n_Body_y[1594] = c_Body_y[1593];
                    end else begin
                        n_Body_x[1594] = c_Body_x[c_Size-1];
                        n_Body_y[1594] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1595) begin
                        n_Body_x[1595] = c_Body_x[1594];
                        n_Body_y[1595] = c_Body_y[1594];
                    end else begin
                        n_Body_x[1595] = c_Body_x[c_Size-1];
                        n_Body_y[1595] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1596) begin
                        n_Body_x[1596] = c_Body_x[1595];
                        n_Body_y[1596] = c_Body_y[1595];
                    end else begin
                        n_Body_x[1596] = c_Body_x[c_Size-1];
                        n_Body_y[1596] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1597) begin
                        n_Body_x[1597] = c_Body_x[1596];
                        n_Body_y[1597] = c_Body_y[1596];
                    end else begin
                        n_Body_x[1597] = c_Body_x[c_Size-1];
                        n_Body_y[1597] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1598) begin
                        n_Body_x[1598] = c_Body_x[1597];
                        n_Body_y[1598] = c_Body_y[1597];
                    end else begin
                        n_Body_x[1598] = c_Body_x[c_Size-1];
                        n_Body_y[1598] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1599) begin
                        n_Body_x[1599] = c_Body_x[1598];
                        n_Body_y[1599] = c_Body_y[1598];
                    end else begin
                        n_Body_x[1599] = c_Body_x[c_Size-1];
                        n_Body_y[1599] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1600) begin
                        n_Body_x[1600] = c_Body_x[1599];
                        n_Body_y[1600] = c_Body_y[1599];
                    end else begin
                        n_Body_x[1600] = c_Body_x[c_Size-1];
                        n_Body_y[1600] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1601) begin
                        n_Body_x[1601] = c_Body_x[1600];
                        n_Body_y[1601] = c_Body_y[1600];
                    end else begin
                        n_Body_x[1601] = c_Body_x[c_Size-1];
                        n_Body_y[1601] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1602) begin
                        n_Body_x[1602] = c_Body_x[1601];
                        n_Body_y[1602] = c_Body_y[1601];
                    end else begin
                        n_Body_x[1602] = c_Body_x[c_Size-1];
                        n_Body_y[1602] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1603) begin
                        n_Body_x[1603] = c_Body_x[1602];
                        n_Body_y[1603] = c_Body_y[1602];
                    end else begin
                        n_Body_x[1603] = c_Body_x[c_Size-1];
                        n_Body_y[1603] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1604) begin
                        n_Body_x[1604] = c_Body_x[1603];
                        n_Body_y[1604] = c_Body_y[1603];
                    end else begin
                        n_Body_x[1604] = c_Body_x[c_Size-1];
                        n_Body_y[1604] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1605) begin
                        n_Body_x[1605] = c_Body_x[1604];
                        n_Body_y[1605] = c_Body_y[1604];
                    end else begin
                        n_Body_x[1605] = c_Body_x[c_Size-1];
                        n_Body_y[1605] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1606) begin
                        n_Body_x[1606] = c_Body_x[1605];
                        n_Body_y[1606] = c_Body_y[1605];
                    end else begin
                        n_Body_x[1606] = c_Body_x[c_Size-1];
                        n_Body_y[1606] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1607) begin
                        n_Body_x[1607] = c_Body_x[1606];
                        n_Body_y[1607] = c_Body_y[1606];
                    end else begin
                        n_Body_x[1607] = c_Body_x[c_Size-1];
                        n_Body_y[1607] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1608) begin
                        n_Body_x[1608] = c_Body_x[1607];
                        n_Body_y[1608] = c_Body_y[1607];
                    end else begin
                        n_Body_x[1608] = c_Body_x[c_Size-1];
                        n_Body_y[1608] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1609) begin
                        n_Body_x[1609] = c_Body_x[1608];
                        n_Body_y[1609] = c_Body_y[1608];
                    end else begin
                        n_Body_x[1609] = c_Body_x[c_Size-1];
                        n_Body_y[1609] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1610) begin
                        n_Body_x[1610] = c_Body_x[1609];
                        n_Body_y[1610] = c_Body_y[1609];
                    end else begin
                        n_Body_x[1610] = c_Body_x[c_Size-1];
                        n_Body_y[1610] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1611) begin
                        n_Body_x[1611] = c_Body_x[1610];
                        n_Body_y[1611] = c_Body_y[1610];
                    end else begin
                        n_Body_x[1611] = c_Body_x[c_Size-1];
                        n_Body_y[1611] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1612) begin
                        n_Body_x[1612] = c_Body_x[1611];
                        n_Body_y[1612] = c_Body_y[1611];
                    end else begin
                        n_Body_x[1612] = c_Body_x[c_Size-1];
                        n_Body_y[1612] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1613) begin
                        n_Body_x[1613] = c_Body_x[1612];
                        n_Body_y[1613] = c_Body_y[1612];
                    end else begin
                        n_Body_x[1613] = c_Body_x[c_Size-1];
                        n_Body_y[1613] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1614) begin
                        n_Body_x[1614] = c_Body_x[1613];
                        n_Body_y[1614] = c_Body_y[1613];
                    end else begin
                        n_Body_x[1614] = c_Body_x[c_Size-1];
                        n_Body_y[1614] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1615) begin
                        n_Body_x[1615] = c_Body_x[1614];
                        n_Body_y[1615] = c_Body_y[1614];
                    end else begin
                        n_Body_x[1615] = c_Body_x[c_Size-1];
                        n_Body_y[1615] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1616) begin
                        n_Body_x[1616] = c_Body_x[1615];
                        n_Body_y[1616] = c_Body_y[1615];
                    end else begin
                        n_Body_x[1616] = c_Body_x[c_Size-1];
                        n_Body_y[1616] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1617) begin
                        n_Body_x[1617] = c_Body_x[1616];
                        n_Body_y[1617] = c_Body_y[1616];
                    end else begin
                        n_Body_x[1617] = c_Body_x[c_Size-1];
                        n_Body_y[1617] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1618) begin
                        n_Body_x[1618] = c_Body_x[1617];
                        n_Body_y[1618] = c_Body_y[1617];
                    end else begin
                        n_Body_x[1618] = c_Body_x[c_Size-1];
                        n_Body_y[1618] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1619) begin
                        n_Body_x[1619] = c_Body_x[1618];
                        n_Body_y[1619] = c_Body_y[1618];
                    end else begin
                        n_Body_x[1619] = c_Body_x[c_Size-1];
                        n_Body_y[1619] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1620) begin
                        n_Body_x[1620] = c_Body_x[1619];
                        n_Body_y[1620] = c_Body_y[1619];
                    end else begin
                        n_Body_x[1620] = c_Body_x[c_Size-1];
                        n_Body_y[1620] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1621) begin
                        n_Body_x[1621] = c_Body_x[1620];
                        n_Body_y[1621] = c_Body_y[1620];
                    end else begin
                        n_Body_x[1621] = c_Body_x[c_Size-1];
                        n_Body_y[1621] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1622) begin
                        n_Body_x[1622] = c_Body_x[1621];
                        n_Body_y[1622] = c_Body_y[1621];
                    end else begin
                        n_Body_x[1622] = c_Body_x[c_Size-1];
                        n_Body_y[1622] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1623) begin
                        n_Body_x[1623] = c_Body_x[1622];
                        n_Body_y[1623] = c_Body_y[1622];
                    end else begin
                        n_Body_x[1623] = c_Body_x[c_Size-1];
                        n_Body_y[1623] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1624) begin
                        n_Body_x[1624] = c_Body_x[1623];
                        n_Body_y[1624] = c_Body_y[1623];
                    end else begin
                        n_Body_x[1624] = c_Body_x[c_Size-1];
                        n_Body_y[1624] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1625) begin
                        n_Body_x[1625] = c_Body_x[1624];
                        n_Body_y[1625] = c_Body_y[1624];
                    end else begin
                        n_Body_x[1625] = c_Body_x[c_Size-1];
                        n_Body_y[1625] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1626) begin
                        n_Body_x[1626] = c_Body_x[1625];
                        n_Body_y[1626] = c_Body_y[1625];
                    end else begin
                        n_Body_x[1626] = c_Body_x[c_Size-1];
                        n_Body_y[1626] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1627) begin
                        n_Body_x[1627] = c_Body_x[1626];
                        n_Body_y[1627] = c_Body_y[1626];
                    end else begin
                        n_Body_x[1627] = c_Body_x[c_Size-1];
                        n_Body_y[1627] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1628) begin
                        n_Body_x[1628] = c_Body_x[1627];
                        n_Body_y[1628] = c_Body_y[1627];
                    end else begin
                        n_Body_x[1628] = c_Body_x[c_Size-1];
                        n_Body_y[1628] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1629) begin
                        n_Body_x[1629] = c_Body_x[1628];
                        n_Body_y[1629] = c_Body_y[1628];
                    end else begin
                        n_Body_x[1629] = c_Body_x[c_Size-1];
                        n_Body_y[1629] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1630) begin
                        n_Body_x[1630] = c_Body_x[1629];
                        n_Body_y[1630] = c_Body_y[1629];
                    end else begin
                        n_Body_x[1630] = c_Body_x[c_Size-1];
                        n_Body_y[1630] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1631) begin
                        n_Body_x[1631] = c_Body_x[1630];
                        n_Body_y[1631] = c_Body_y[1630];
                    end else begin
                        n_Body_x[1631] = c_Body_x[c_Size-1];
                        n_Body_y[1631] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1632) begin
                        n_Body_x[1632] = c_Body_x[1631];
                        n_Body_y[1632] = c_Body_y[1631];
                    end else begin
                        n_Body_x[1632] = c_Body_x[c_Size-1];
                        n_Body_y[1632] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1633) begin
                        n_Body_x[1633] = c_Body_x[1632];
                        n_Body_y[1633] = c_Body_y[1632];
                    end else begin
                        n_Body_x[1633] = c_Body_x[c_Size-1];
                        n_Body_y[1633] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1634) begin
                        n_Body_x[1634] = c_Body_x[1633];
                        n_Body_y[1634] = c_Body_y[1633];
                    end else begin
                        n_Body_x[1634] = c_Body_x[c_Size-1];
                        n_Body_y[1634] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1635) begin
                        n_Body_x[1635] = c_Body_x[1634];
                        n_Body_y[1635] = c_Body_y[1634];
                    end else begin
                        n_Body_x[1635] = c_Body_x[c_Size-1];
                        n_Body_y[1635] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1636) begin
                        n_Body_x[1636] = c_Body_x[1635];
                        n_Body_y[1636] = c_Body_y[1635];
                    end else begin
                        n_Body_x[1636] = c_Body_x[c_Size-1];
                        n_Body_y[1636] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1637) begin
                        n_Body_x[1637] = c_Body_x[1636];
                        n_Body_y[1637] = c_Body_y[1636];
                    end else begin
                        n_Body_x[1637] = c_Body_x[c_Size-1];
                        n_Body_y[1637] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1638) begin
                        n_Body_x[1638] = c_Body_x[1637];
                        n_Body_y[1638] = c_Body_y[1637];
                    end else begin
                        n_Body_x[1638] = c_Body_x[c_Size-1];
                        n_Body_y[1638] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1639) begin
                        n_Body_x[1639] = c_Body_x[1638];
                        n_Body_y[1639] = c_Body_y[1638];
                    end else begin
                        n_Body_x[1639] = c_Body_x[c_Size-1];
                        n_Body_y[1639] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1640) begin
                        n_Body_x[1640] = c_Body_x[1639];
                        n_Body_y[1640] = c_Body_y[1639];
                    end else begin
                        n_Body_x[1640] = c_Body_x[c_Size-1];
                        n_Body_y[1640] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1641) begin
                        n_Body_x[1641] = c_Body_x[1640];
                        n_Body_y[1641] = c_Body_y[1640];
                    end else begin
                        n_Body_x[1641] = c_Body_x[c_Size-1];
                        n_Body_y[1641] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1642) begin
                        n_Body_x[1642] = c_Body_x[1641];
                        n_Body_y[1642] = c_Body_y[1641];
                    end else begin
                        n_Body_x[1642] = c_Body_x[c_Size-1];
                        n_Body_y[1642] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1643) begin
                        n_Body_x[1643] = c_Body_x[1642];
                        n_Body_y[1643] = c_Body_y[1642];
                    end else begin
                        n_Body_x[1643] = c_Body_x[c_Size-1];
                        n_Body_y[1643] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1644) begin
                        n_Body_x[1644] = c_Body_x[1643];
                        n_Body_y[1644] = c_Body_y[1643];
                    end else begin
                        n_Body_x[1644] = c_Body_x[c_Size-1];
                        n_Body_y[1644] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1645) begin
                        n_Body_x[1645] = c_Body_x[1644];
                        n_Body_y[1645] = c_Body_y[1644];
                    end else begin
                        n_Body_x[1645] = c_Body_x[c_Size-1];
                        n_Body_y[1645] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1646) begin
                        n_Body_x[1646] = c_Body_x[1645];
                        n_Body_y[1646] = c_Body_y[1645];
                    end else begin
                        n_Body_x[1646] = c_Body_x[c_Size-1];
                        n_Body_y[1646] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1647) begin
                        n_Body_x[1647] = c_Body_x[1646];
                        n_Body_y[1647] = c_Body_y[1646];
                    end else begin
                        n_Body_x[1647] = c_Body_x[c_Size-1];
                        n_Body_y[1647] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1648) begin
                        n_Body_x[1648] = c_Body_x[1647];
                        n_Body_y[1648] = c_Body_y[1647];
                    end else begin
                        n_Body_x[1648] = c_Body_x[c_Size-1];
                        n_Body_y[1648] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1649) begin
                        n_Body_x[1649] = c_Body_x[1648];
                        n_Body_y[1649] = c_Body_y[1648];
                    end else begin
                        n_Body_x[1649] = c_Body_x[c_Size-1];
                        n_Body_y[1649] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1650) begin
                        n_Body_x[1650] = c_Body_x[1649];
                        n_Body_y[1650] = c_Body_y[1649];
                    end else begin
                        n_Body_x[1650] = c_Body_x[c_Size-1];
                        n_Body_y[1650] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1651) begin
                        n_Body_x[1651] = c_Body_x[1650];
                        n_Body_y[1651] = c_Body_y[1650];
                    end else begin
                        n_Body_x[1651] = c_Body_x[c_Size-1];
                        n_Body_y[1651] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1652) begin
                        n_Body_x[1652] = c_Body_x[1651];
                        n_Body_y[1652] = c_Body_y[1651];
                    end else begin
                        n_Body_x[1652] = c_Body_x[c_Size-1];
                        n_Body_y[1652] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1653) begin
                        n_Body_x[1653] = c_Body_x[1652];
                        n_Body_y[1653] = c_Body_y[1652];
                    end else begin
                        n_Body_x[1653] = c_Body_x[c_Size-1];
                        n_Body_y[1653] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1654) begin
                        n_Body_x[1654] = c_Body_x[1653];
                        n_Body_y[1654] = c_Body_y[1653];
                    end else begin
                        n_Body_x[1654] = c_Body_x[c_Size-1];
                        n_Body_y[1654] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1655) begin
                        n_Body_x[1655] = c_Body_x[1654];
                        n_Body_y[1655] = c_Body_y[1654];
                    end else begin
                        n_Body_x[1655] = c_Body_x[c_Size-1];
                        n_Body_y[1655] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1656) begin
                        n_Body_x[1656] = c_Body_x[1655];
                        n_Body_y[1656] = c_Body_y[1655];
                    end else begin
                        n_Body_x[1656] = c_Body_x[c_Size-1];
                        n_Body_y[1656] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1657) begin
                        n_Body_x[1657] = c_Body_x[1656];
                        n_Body_y[1657] = c_Body_y[1656];
                    end else begin
                        n_Body_x[1657] = c_Body_x[c_Size-1];
                        n_Body_y[1657] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1658) begin
                        n_Body_x[1658] = c_Body_x[1657];
                        n_Body_y[1658] = c_Body_y[1657];
                    end else begin
                        n_Body_x[1658] = c_Body_x[c_Size-1];
                        n_Body_y[1658] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1659) begin
                        n_Body_x[1659] = c_Body_x[1658];
                        n_Body_y[1659] = c_Body_y[1658];
                    end else begin
                        n_Body_x[1659] = c_Body_x[c_Size-1];
                        n_Body_y[1659] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1660) begin
                        n_Body_x[1660] = c_Body_x[1659];
                        n_Body_y[1660] = c_Body_y[1659];
                    end else begin
                        n_Body_x[1660] = c_Body_x[c_Size-1];
                        n_Body_y[1660] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1661) begin
                        n_Body_x[1661] = c_Body_x[1660];
                        n_Body_y[1661] = c_Body_y[1660];
                    end else begin
                        n_Body_x[1661] = c_Body_x[c_Size-1];
                        n_Body_y[1661] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1662) begin
                        n_Body_x[1662] = c_Body_x[1661];
                        n_Body_y[1662] = c_Body_y[1661];
                    end else begin
                        n_Body_x[1662] = c_Body_x[c_Size-1];
                        n_Body_y[1662] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1663) begin
                        n_Body_x[1663] = c_Body_x[1662];
                        n_Body_y[1663] = c_Body_y[1662];
                    end else begin
                        n_Body_x[1663] = c_Body_x[c_Size-1];
                        n_Body_y[1663] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1664) begin
                        n_Body_x[1664] = c_Body_x[1663];
                        n_Body_y[1664] = c_Body_y[1663];
                    end else begin
                        n_Body_x[1664] = c_Body_x[c_Size-1];
                        n_Body_y[1664] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1665) begin
                        n_Body_x[1665] = c_Body_x[1664];
                        n_Body_y[1665] = c_Body_y[1664];
                    end else begin
                        n_Body_x[1665] = c_Body_x[c_Size-1];
                        n_Body_y[1665] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1666) begin
                        n_Body_x[1666] = c_Body_x[1665];
                        n_Body_y[1666] = c_Body_y[1665];
                    end else begin
                        n_Body_x[1666] = c_Body_x[c_Size-1];
                        n_Body_y[1666] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1667) begin
                        n_Body_x[1667] = c_Body_x[1666];
                        n_Body_y[1667] = c_Body_y[1666];
                    end else begin
                        n_Body_x[1667] = c_Body_x[c_Size-1];
                        n_Body_y[1667] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1668) begin
                        n_Body_x[1668] = c_Body_x[1667];
                        n_Body_y[1668] = c_Body_y[1667];
                    end else begin
                        n_Body_x[1668] = c_Body_x[c_Size-1];
                        n_Body_y[1668] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1669) begin
                        n_Body_x[1669] = c_Body_x[1668];
                        n_Body_y[1669] = c_Body_y[1668];
                    end else begin
                        n_Body_x[1669] = c_Body_x[c_Size-1];
                        n_Body_y[1669] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1670) begin
                        n_Body_x[1670] = c_Body_x[1669];
                        n_Body_y[1670] = c_Body_y[1669];
                    end else begin
                        n_Body_x[1670] = c_Body_x[c_Size-1];
                        n_Body_y[1670] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1671) begin
                        n_Body_x[1671] = c_Body_x[1670];
                        n_Body_y[1671] = c_Body_y[1670];
                    end else begin
                        n_Body_x[1671] = c_Body_x[c_Size-1];
                        n_Body_y[1671] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1672) begin
                        n_Body_x[1672] = c_Body_x[1671];
                        n_Body_y[1672] = c_Body_y[1671];
                    end else begin
                        n_Body_x[1672] = c_Body_x[c_Size-1];
                        n_Body_y[1672] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1673) begin
                        n_Body_x[1673] = c_Body_x[1672];
                        n_Body_y[1673] = c_Body_y[1672];
                    end else begin
                        n_Body_x[1673] = c_Body_x[c_Size-1];
                        n_Body_y[1673] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1674) begin
                        n_Body_x[1674] = c_Body_x[1673];
                        n_Body_y[1674] = c_Body_y[1673];
                    end else begin
                        n_Body_x[1674] = c_Body_x[c_Size-1];
                        n_Body_y[1674] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1675) begin
                        n_Body_x[1675] = c_Body_x[1674];
                        n_Body_y[1675] = c_Body_y[1674];
                    end else begin
                        n_Body_x[1675] = c_Body_x[c_Size-1];
                        n_Body_y[1675] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1676) begin
                        n_Body_x[1676] = c_Body_x[1675];
                        n_Body_y[1676] = c_Body_y[1675];
                    end else begin
                        n_Body_x[1676] = c_Body_x[c_Size-1];
                        n_Body_y[1676] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1677) begin
                        n_Body_x[1677] = c_Body_x[1676];
                        n_Body_y[1677] = c_Body_y[1676];
                    end else begin
                        n_Body_x[1677] = c_Body_x[c_Size-1];
                        n_Body_y[1677] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1678) begin
                        n_Body_x[1678] = c_Body_x[1677];
                        n_Body_y[1678] = c_Body_y[1677];
                    end else begin
                        n_Body_x[1678] = c_Body_x[c_Size-1];
                        n_Body_y[1678] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1679) begin
                        n_Body_x[1679] = c_Body_x[1678];
                        n_Body_y[1679] = c_Body_y[1678];
                    end else begin
                        n_Body_x[1679] = c_Body_x[c_Size-1];
                        n_Body_y[1679] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1680) begin
                        n_Body_x[1680] = c_Body_x[1679];
                        n_Body_y[1680] = c_Body_y[1679];
                    end else begin
                        n_Body_x[1680] = c_Body_x[c_Size-1];
                        n_Body_y[1680] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1681) begin
                        n_Body_x[1681] = c_Body_x[1680];
                        n_Body_y[1681] = c_Body_y[1680];
                    end else begin
                        n_Body_x[1681] = c_Body_x[c_Size-1];
                        n_Body_y[1681] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1682) begin
                        n_Body_x[1682] = c_Body_x[1681];
                        n_Body_y[1682] = c_Body_y[1681];
                    end else begin
                        n_Body_x[1682] = c_Body_x[c_Size-1];
                        n_Body_y[1682] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1683) begin
                        n_Body_x[1683] = c_Body_x[1682];
                        n_Body_y[1683] = c_Body_y[1682];
                    end else begin
                        n_Body_x[1683] = c_Body_x[c_Size-1];
                        n_Body_y[1683] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1684) begin
                        n_Body_x[1684] = c_Body_x[1683];
                        n_Body_y[1684] = c_Body_y[1683];
                    end else begin
                        n_Body_x[1684] = c_Body_x[c_Size-1];
                        n_Body_y[1684] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1685) begin
                        n_Body_x[1685] = c_Body_x[1684];
                        n_Body_y[1685] = c_Body_y[1684];
                    end else begin
                        n_Body_x[1685] = c_Body_x[c_Size-1];
                        n_Body_y[1685] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1686) begin
                        n_Body_x[1686] = c_Body_x[1685];
                        n_Body_y[1686] = c_Body_y[1685];
                    end else begin
                        n_Body_x[1686] = c_Body_x[c_Size-1];
                        n_Body_y[1686] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1687) begin
                        n_Body_x[1687] = c_Body_x[1686];
                        n_Body_y[1687] = c_Body_y[1686];
                    end else begin
                        n_Body_x[1687] = c_Body_x[c_Size-1];
                        n_Body_y[1687] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1688) begin
                        n_Body_x[1688] = c_Body_x[1687];
                        n_Body_y[1688] = c_Body_y[1687];
                    end else begin
                        n_Body_x[1688] = c_Body_x[c_Size-1];
                        n_Body_y[1688] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1689) begin
                        n_Body_x[1689] = c_Body_x[1688];
                        n_Body_y[1689] = c_Body_y[1688];
                    end else begin
                        n_Body_x[1689] = c_Body_x[c_Size-1];
                        n_Body_y[1689] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1690) begin
                        n_Body_x[1690] = c_Body_x[1689];
                        n_Body_y[1690] = c_Body_y[1689];
                    end else begin
                        n_Body_x[1690] = c_Body_x[c_Size-1];
                        n_Body_y[1690] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1691) begin
                        n_Body_x[1691] = c_Body_x[1690];
                        n_Body_y[1691] = c_Body_y[1690];
                    end else begin
                        n_Body_x[1691] = c_Body_x[c_Size-1];
                        n_Body_y[1691] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1692) begin
                        n_Body_x[1692] = c_Body_x[1691];
                        n_Body_y[1692] = c_Body_y[1691];
                    end else begin
                        n_Body_x[1692] = c_Body_x[c_Size-1];
                        n_Body_y[1692] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1693) begin
                        n_Body_x[1693] = c_Body_x[1692];
                        n_Body_y[1693] = c_Body_y[1692];
                    end else begin
                        n_Body_x[1693] = c_Body_x[c_Size-1];
                        n_Body_y[1693] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1694) begin
                        n_Body_x[1694] = c_Body_x[1693];
                        n_Body_y[1694] = c_Body_y[1693];
                    end else begin
                        n_Body_x[1694] = c_Body_x[c_Size-1];
                        n_Body_y[1694] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1695) begin
                        n_Body_x[1695] = c_Body_x[1694];
                        n_Body_y[1695] = c_Body_y[1694];
                    end else begin
                        n_Body_x[1695] = c_Body_x[c_Size-1];
                        n_Body_y[1695] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1696) begin
                        n_Body_x[1696] = c_Body_x[1695];
                        n_Body_y[1696] = c_Body_y[1695];
                    end else begin
                        n_Body_x[1696] = c_Body_x[c_Size-1];
                        n_Body_y[1696] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1697) begin
                        n_Body_x[1697] = c_Body_x[1696];
                        n_Body_y[1697] = c_Body_y[1696];
                    end else begin
                        n_Body_x[1697] = c_Body_x[c_Size-1];
                        n_Body_y[1697] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1698) begin
                        n_Body_x[1698] = c_Body_x[1697];
                        n_Body_y[1698] = c_Body_y[1697];
                    end else begin
                        n_Body_x[1698] = c_Body_x[c_Size-1];
                        n_Body_y[1698] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1699) begin
                        n_Body_x[1699] = c_Body_x[1698];
                        n_Body_y[1699] = c_Body_y[1698];
                    end else begin
                        n_Body_x[1699] = c_Body_x[c_Size-1];
                        n_Body_y[1699] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1700) begin
                        n_Body_x[1700] = c_Body_x[1699];
                        n_Body_y[1700] = c_Body_y[1699];
                    end else begin
                        n_Body_x[1700] = c_Body_x[c_Size-1];
                        n_Body_y[1700] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1701) begin
                        n_Body_x[1701] = c_Body_x[1700];
                        n_Body_y[1701] = c_Body_y[1700];
                    end else begin
                        n_Body_x[1701] = c_Body_x[c_Size-1];
                        n_Body_y[1701] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1702) begin
                        n_Body_x[1702] = c_Body_x[1701];
                        n_Body_y[1702] = c_Body_y[1701];
                    end else begin
                        n_Body_x[1702] = c_Body_x[c_Size-1];
                        n_Body_y[1702] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1703) begin
                        n_Body_x[1703] = c_Body_x[1702];
                        n_Body_y[1703] = c_Body_y[1702];
                    end else begin
                        n_Body_x[1703] = c_Body_x[c_Size-1];
                        n_Body_y[1703] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1704) begin
                        n_Body_x[1704] = c_Body_x[1703];
                        n_Body_y[1704] = c_Body_y[1703];
                    end else begin
                        n_Body_x[1704] = c_Body_x[c_Size-1];
                        n_Body_y[1704] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1705) begin
                        n_Body_x[1705] = c_Body_x[1704];
                        n_Body_y[1705] = c_Body_y[1704];
                    end else begin
                        n_Body_x[1705] = c_Body_x[c_Size-1];
                        n_Body_y[1705] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1706) begin
                        n_Body_x[1706] = c_Body_x[1705];
                        n_Body_y[1706] = c_Body_y[1705];
                    end else begin
                        n_Body_x[1706] = c_Body_x[c_Size-1];
                        n_Body_y[1706] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1707) begin
                        n_Body_x[1707] = c_Body_x[1706];
                        n_Body_y[1707] = c_Body_y[1706];
                    end else begin
                        n_Body_x[1707] = c_Body_x[c_Size-1];
                        n_Body_y[1707] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1708) begin
                        n_Body_x[1708] = c_Body_x[1707];
                        n_Body_y[1708] = c_Body_y[1707];
                    end else begin
                        n_Body_x[1708] = c_Body_x[c_Size-1];
                        n_Body_y[1708] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1709) begin
                        n_Body_x[1709] = c_Body_x[1708];
                        n_Body_y[1709] = c_Body_y[1708];
                    end else begin
                        n_Body_x[1709] = c_Body_x[c_Size-1];
                        n_Body_y[1709] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1710) begin
                        n_Body_x[1710] = c_Body_x[1709];
                        n_Body_y[1710] = c_Body_y[1709];
                    end else begin
                        n_Body_x[1710] = c_Body_x[c_Size-1];
                        n_Body_y[1710] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1711) begin
                        n_Body_x[1711] = c_Body_x[1710];
                        n_Body_y[1711] = c_Body_y[1710];
                    end else begin
                        n_Body_x[1711] = c_Body_x[c_Size-1];
                        n_Body_y[1711] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1712) begin
                        n_Body_x[1712] = c_Body_x[1711];
                        n_Body_y[1712] = c_Body_y[1711];
                    end else begin
                        n_Body_x[1712] = c_Body_x[c_Size-1];
                        n_Body_y[1712] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1713) begin
                        n_Body_x[1713] = c_Body_x[1712];
                        n_Body_y[1713] = c_Body_y[1712];
                    end else begin
                        n_Body_x[1713] = c_Body_x[c_Size-1];
                        n_Body_y[1713] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1714) begin
                        n_Body_x[1714] = c_Body_x[1713];
                        n_Body_y[1714] = c_Body_y[1713];
                    end else begin
                        n_Body_x[1714] = c_Body_x[c_Size-1];
                        n_Body_y[1714] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1715) begin
                        n_Body_x[1715] = c_Body_x[1714];
                        n_Body_y[1715] = c_Body_y[1714];
                    end else begin
                        n_Body_x[1715] = c_Body_x[c_Size-1];
                        n_Body_y[1715] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1716) begin
                        n_Body_x[1716] = c_Body_x[1715];
                        n_Body_y[1716] = c_Body_y[1715];
                    end else begin
                        n_Body_x[1716] = c_Body_x[c_Size-1];
                        n_Body_y[1716] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1717) begin
                        n_Body_x[1717] = c_Body_x[1716];
                        n_Body_y[1717] = c_Body_y[1716];
                    end else begin
                        n_Body_x[1717] = c_Body_x[c_Size-1];
                        n_Body_y[1717] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1718) begin
                        n_Body_x[1718] = c_Body_x[1717];
                        n_Body_y[1718] = c_Body_y[1717];
                    end else begin
                        n_Body_x[1718] = c_Body_x[c_Size-1];
                        n_Body_y[1718] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1719) begin
                        n_Body_x[1719] = c_Body_x[1718];
                        n_Body_y[1719] = c_Body_y[1718];
                    end else begin
                        n_Body_x[1719] = c_Body_x[c_Size-1];
                        n_Body_y[1719] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1720) begin
                        n_Body_x[1720] = c_Body_x[1719];
                        n_Body_y[1720] = c_Body_y[1719];
                    end else begin
                        n_Body_x[1720] = c_Body_x[c_Size-1];
                        n_Body_y[1720] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1721) begin
                        n_Body_x[1721] = c_Body_x[1720];
                        n_Body_y[1721] = c_Body_y[1720];
                    end else begin
                        n_Body_x[1721] = c_Body_x[c_Size-1];
                        n_Body_y[1721] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1722) begin
                        n_Body_x[1722] = c_Body_x[1721];
                        n_Body_y[1722] = c_Body_y[1721];
                    end else begin
                        n_Body_x[1722] = c_Body_x[c_Size-1];
                        n_Body_y[1722] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1723) begin
                        n_Body_x[1723] = c_Body_x[1722];
                        n_Body_y[1723] = c_Body_y[1722];
                    end else begin
                        n_Body_x[1723] = c_Body_x[c_Size-1];
                        n_Body_y[1723] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1724) begin
                        n_Body_x[1724] = c_Body_x[1723];
                        n_Body_y[1724] = c_Body_y[1723];
                    end else begin
                        n_Body_x[1724] = c_Body_x[c_Size-1];
                        n_Body_y[1724] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1725) begin
                        n_Body_x[1725] = c_Body_x[1724];
                        n_Body_y[1725] = c_Body_y[1724];
                    end else begin
                        n_Body_x[1725] = c_Body_x[c_Size-1];
                        n_Body_y[1725] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1726) begin
                        n_Body_x[1726] = c_Body_x[1725];
                        n_Body_y[1726] = c_Body_y[1725];
                    end else begin
                        n_Body_x[1726] = c_Body_x[c_Size-1];
                        n_Body_y[1726] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1727) begin
                        n_Body_x[1727] = c_Body_x[1726];
                        n_Body_y[1727] = c_Body_y[1726];
                    end else begin
                        n_Body_x[1727] = c_Body_x[c_Size-1];
                        n_Body_y[1727] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1728) begin
                        n_Body_x[1728] = c_Body_x[1727];
                        n_Body_y[1728] = c_Body_y[1727];
                    end else begin
                        n_Body_x[1728] = c_Body_x[c_Size-1];
                        n_Body_y[1728] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1729) begin
                        n_Body_x[1729] = c_Body_x[1728];
                        n_Body_y[1729] = c_Body_y[1728];
                    end else begin
                        n_Body_x[1729] = c_Body_x[c_Size-1];
                        n_Body_y[1729] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1730) begin
                        n_Body_x[1730] = c_Body_x[1729];
                        n_Body_y[1730] = c_Body_y[1729];
                    end else begin
                        n_Body_x[1730] = c_Body_x[c_Size-1];
                        n_Body_y[1730] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1731) begin
                        n_Body_x[1731] = c_Body_x[1730];
                        n_Body_y[1731] = c_Body_y[1730];
                    end else begin
                        n_Body_x[1731] = c_Body_x[c_Size-1];
                        n_Body_y[1731] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1732) begin
                        n_Body_x[1732] = c_Body_x[1731];
                        n_Body_y[1732] = c_Body_y[1731];
                    end else begin
                        n_Body_x[1732] = c_Body_x[c_Size-1];
                        n_Body_y[1732] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1733) begin
                        n_Body_x[1733] = c_Body_x[1732];
                        n_Body_y[1733] = c_Body_y[1732];
                    end else begin
                        n_Body_x[1733] = c_Body_x[c_Size-1];
                        n_Body_y[1733] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1734) begin
                        n_Body_x[1734] = c_Body_x[1733];
                        n_Body_y[1734] = c_Body_y[1733];
                    end else begin
                        n_Body_x[1734] = c_Body_x[c_Size-1];
                        n_Body_y[1734] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1735) begin
                        n_Body_x[1735] = c_Body_x[1734];
                        n_Body_y[1735] = c_Body_y[1734];
                    end else begin
                        n_Body_x[1735] = c_Body_x[c_Size-1];
                        n_Body_y[1735] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1736) begin
                        n_Body_x[1736] = c_Body_x[1735];
                        n_Body_y[1736] = c_Body_y[1735];
                    end else begin
                        n_Body_x[1736] = c_Body_x[c_Size-1];
                        n_Body_y[1736] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1737) begin
                        n_Body_x[1737] = c_Body_x[1736];
                        n_Body_y[1737] = c_Body_y[1736];
                    end else begin
                        n_Body_x[1737] = c_Body_x[c_Size-1];
                        n_Body_y[1737] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1738) begin
                        n_Body_x[1738] = c_Body_x[1737];
                        n_Body_y[1738] = c_Body_y[1737];
                    end else begin
                        n_Body_x[1738] = c_Body_x[c_Size-1];
                        n_Body_y[1738] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1739) begin
                        n_Body_x[1739] = c_Body_x[1738];
                        n_Body_y[1739] = c_Body_y[1738];
                    end else begin
                        n_Body_x[1739] = c_Body_x[c_Size-1];
                        n_Body_y[1739] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1740) begin
                        n_Body_x[1740] = c_Body_x[1739];
                        n_Body_y[1740] = c_Body_y[1739];
                    end else begin
                        n_Body_x[1740] = c_Body_x[c_Size-1];
                        n_Body_y[1740] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1741) begin
                        n_Body_x[1741] = c_Body_x[1740];
                        n_Body_y[1741] = c_Body_y[1740];
                    end else begin
                        n_Body_x[1741] = c_Body_x[c_Size-1];
                        n_Body_y[1741] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1742) begin
                        n_Body_x[1742] = c_Body_x[1741];
                        n_Body_y[1742] = c_Body_y[1741];
                    end else begin
                        n_Body_x[1742] = c_Body_x[c_Size-1];
                        n_Body_y[1742] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1743) begin
                        n_Body_x[1743] = c_Body_x[1742];
                        n_Body_y[1743] = c_Body_y[1742];
                    end else begin
                        n_Body_x[1743] = c_Body_x[c_Size-1];
                        n_Body_y[1743] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1744) begin
                        n_Body_x[1744] = c_Body_x[1743];
                        n_Body_y[1744] = c_Body_y[1743];
                    end else begin
                        n_Body_x[1744] = c_Body_x[c_Size-1];
                        n_Body_y[1744] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1745) begin
                        n_Body_x[1745] = c_Body_x[1744];
                        n_Body_y[1745] = c_Body_y[1744];
                    end else begin
                        n_Body_x[1745] = c_Body_x[c_Size-1];
                        n_Body_y[1745] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1746) begin
                        n_Body_x[1746] = c_Body_x[1745];
                        n_Body_y[1746] = c_Body_y[1745];
                    end else begin
                        n_Body_x[1746] = c_Body_x[c_Size-1];
                        n_Body_y[1746] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1747) begin
                        n_Body_x[1747] = c_Body_x[1746];
                        n_Body_y[1747] = c_Body_y[1746];
                    end else begin
                        n_Body_x[1747] = c_Body_x[c_Size-1];
                        n_Body_y[1747] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1748) begin
                        n_Body_x[1748] = c_Body_x[1747];
                        n_Body_y[1748] = c_Body_y[1747];
                    end else begin
                        n_Body_x[1748] = c_Body_x[c_Size-1];
                        n_Body_y[1748] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1749) begin
                        n_Body_x[1749] = c_Body_x[1748];
                        n_Body_y[1749] = c_Body_y[1748];
                    end else begin
                        n_Body_x[1749] = c_Body_x[c_Size-1];
                        n_Body_y[1749] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1750) begin
                        n_Body_x[1750] = c_Body_x[1749];
                        n_Body_y[1750] = c_Body_y[1749];
                    end else begin
                        n_Body_x[1750] = c_Body_x[c_Size-1];
                        n_Body_y[1750] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1751) begin
                        n_Body_x[1751] = c_Body_x[1750];
                        n_Body_y[1751] = c_Body_y[1750];
                    end else begin
                        n_Body_x[1751] = c_Body_x[c_Size-1];
                        n_Body_y[1751] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1752) begin
                        n_Body_x[1752] = c_Body_x[1751];
                        n_Body_y[1752] = c_Body_y[1751];
                    end else begin
                        n_Body_x[1752] = c_Body_x[c_Size-1];
                        n_Body_y[1752] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1753) begin
                        n_Body_x[1753] = c_Body_x[1752];
                        n_Body_y[1753] = c_Body_y[1752];
                    end else begin
                        n_Body_x[1753] = c_Body_x[c_Size-1];
                        n_Body_y[1753] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1754) begin
                        n_Body_x[1754] = c_Body_x[1753];
                        n_Body_y[1754] = c_Body_y[1753];
                    end else begin
                        n_Body_x[1754] = c_Body_x[c_Size-1];
                        n_Body_y[1754] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1755) begin
                        n_Body_x[1755] = c_Body_x[1754];
                        n_Body_y[1755] = c_Body_y[1754];
                    end else begin
                        n_Body_x[1755] = c_Body_x[c_Size-1];
                        n_Body_y[1755] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1756) begin
                        n_Body_x[1756] = c_Body_x[1755];
                        n_Body_y[1756] = c_Body_y[1755];
                    end else begin
                        n_Body_x[1756] = c_Body_x[c_Size-1];
                        n_Body_y[1756] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1757) begin
                        n_Body_x[1757] = c_Body_x[1756];
                        n_Body_y[1757] = c_Body_y[1756];
                    end else begin
                        n_Body_x[1757] = c_Body_x[c_Size-1];
                        n_Body_y[1757] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1758) begin
                        n_Body_x[1758] = c_Body_x[1757];
                        n_Body_y[1758] = c_Body_y[1757];
                    end else begin
                        n_Body_x[1758] = c_Body_x[c_Size-1];
                        n_Body_y[1758] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1759) begin
                        n_Body_x[1759] = c_Body_x[1758];
                        n_Body_y[1759] = c_Body_y[1758];
                    end else begin
                        n_Body_x[1759] = c_Body_x[c_Size-1];
                        n_Body_y[1759] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1760) begin
                        n_Body_x[1760] = c_Body_x[1759];
                        n_Body_y[1760] = c_Body_y[1759];
                    end else begin
                        n_Body_x[1760] = c_Body_x[c_Size-1];
                        n_Body_y[1760] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1761) begin
                        n_Body_x[1761] = c_Body_x[1760];
                        n_Body_y[1761] = c_Body_y[1760];
                    end else begin
                        n_Body_x[1761] = c_Body_x[c_Size-1];
                        n_Body_y[1761] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1762) begin
                        n_Body_x[1762] = c_Body_x[1761];
                        n_Body_y[1762] = c_Body_y[1761];
                    end else begin
                        n_Body_x[1762] = c_Body_x[c_Size-1];
                        n_Body_y[1762] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1763) begin
                        n_Body_x[1763] = c_Body_x[1762];
                        n_Body_y[1763] = c_Body_y[1762];
                    end else begin
                        n_Body_x[1763] = c_Body_x[c_Size-1];
                        n_Body_y[1763] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1764) begin
                        n_Body_x[1764] = c_Body_x[1763];
                        n_Body_y[1764] = c_Body_y[1763];
                    end else begin
                        n_Body_x[1764] = c_Body_x[c_Size-1];
                        n_Body_y[1764] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1765) begin
                        n_Body_x[1765] = c_Body_x[1764];
                        n_Body_y[1765] = c_Body_y[1764];
                    end else begin
                        n_Body_x[1765] = c_Body_x[c_Size-1];
                        n_Body_y[1765] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1766) begin
                        n_Body_x[1766] = c_Body_x[1765];
                        n_Body_y[1766] = c_Body_y[1765];
                    end else begin
                        n_Body_x[1766] = c_Body_x[c_Size-1];
                        n_Body_y[1766] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1767) begin
                        n_Body_x[1767] = c_Body_x[1766];
                        n_Body_y[1767] = c_Body_y[1766];
                    end else begin
                        n_Body_x[1767] = c_Body_x[c_Size-1];
                        n_Body_y[1767] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1768) begin
                        n_Body_x[1768] = c_Body_x[1767];
                        n_Body_y[1768] = c_Body_y[1767];
                    end else begin
                        n_Body_x[1768] = c_Body_x[c_Size-1];
                        n_Body_y[1768] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1769) begin
                        n_Body_x[1769] = c_Body_x[1768];
                        n_Body_y[1769] = c_Body_y[1768];
                    end else begin
                        n_Body_x[1769] = c_Body_x[c_Size-1];
                        n_Body_y[1769] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1770) begin
                        n_Body_x[1770] = c_Body_x[1769];
                        n_Body_y[1770] = c_Body_y[1769];
                    end else begin
                        n_Body_x[1770] = c_Body_x[c_Size-1];
                        n_Body_y[1770] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1771) begin
                        n_Body_x[1771] = c_Body_x[1770];
                        n_Body_y[1771] = c_Body_y[1770];
                    end else begin
                        n_Body_x[1771] = c_Body_x[c_Size-1];
                        n_Body_y[1771] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1772) begin
                        n_Body_x[1772] = c_Body_x[1771];
                        n_Body_y[1772] = c_Body_y[1771];
                    end else begin
                        n_Body_x[1772] = c_Body_x[c_Size-1];
                        n_Body_y[1772] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1773) begin
                        n_Body_x[1773] = c_Body_x[1772];
                        n_Body_y[1773] = c_Body_y[1772];
                    end else begin
                        n_Body_x[1773] = c_Body_x[c_Size-1];
                        n_Body_y[1773] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1774) begin
                        n_Body_x[1774] = c_Body_x[1773];
                        n_Body_y[1774] = c_Body_y[1773];
                    end else begin
                        n_Body_x[1774] = c_Body_x[c_Size-1];
                        n_Body_y[1774] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1775) begin
                        n_Body_x[1775] = c_Body_x[1774];
                        n_Body_y[1775] = c_Body_y[1774];
                    end else begin
                        n_Body_x[1775] = c_Body_x[c_Size-1];
                        n_Body_y[1775] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1776) begin
                        n_Body_x[1776] = c_Body_x[1775];
                        n_Body_y[1776] = c_Body_y[1775];
                    end else begin
                        n_Body_x[1776] = c_Body_x[c_Size-1];
                        n_Body_y[1776] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1777) begin
                        n_Body_x[1777] = c_Body_x[1776];
                        n_Body_y[1777] = c_Body_y[1776];
                    end else begin
                        n_Body_x[1777] = c_Body_x[c_Size-1];
                        n_Body_y[1777] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1778) begin
                        n_Body_x[1778] = c_Body_x[1777];
                        n_Body_y[1778] = c_Body_y[1777];
                    end else begin
                        n_Body_x[1778] = c_Body_x[c_Size-1];
                        n_Body_y[1778] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1779) begin
                        n_Body_x[1779] = c_Body_x[1778];
                        n_Body_y[1779] = c_Body_y[1778];
                    end else begin
                        n_Body_x[1779] = c_Body_x[c_Size-1];
                        n_Body_y[1779] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1780) begin
                        n_Body_x[1780] = c_Body_x[1779];
                        n_Body_y[1780] = c_Body_y[1779];
                    end else begin
                        n_Body_x[1780] = c_Body_x[c_Size-1];
                        n_Body_y[1780] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1781) begin
                        n_Body_x[1781] = c_Body_x[1780];
                        n_Body_y[1781] = c_Body_y[1780];
                    end else begin
                        n_Body_x[1781] = c_Body_x[c_Size-1];
                        n_Body_y[1781] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1782) begin
                        n_Body_x[1782] = c_Body_x[1781];
                        n_Body_y[1782] = c_Body_y[1781];
                    end else begin
                        n_Body_x[1782] = c_Body_x[c_Size-1];
                        n_Body_y[1782] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1783) begin
                        n_Body_x[1783] = c_Body_x[1782];
                        n_Body_y[1783] = c_Body_y[1782];
                    end else begin
                        n_Body_x[1783] = c_Body_x[c_Size-1];
                        n_Body_y[1783] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1784) begin
                        n_Body_x[1784] = c_Body_x[1783];
                        n_Body_y[1784] = c_Body_y[1783];
                    end else begin
                        n_Body_x[1784] = c_Body_x[c_Size-1];
                        n_Body_y[1784] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1785) begin
                        n_Body_x[1785] = c_Body_x[1784];
                        n_Body_y[1785] = c_Body_y[1784];
                    end else begin
                        n_Body_x[1785] = c_Body_x[c_Size-1];
                        n_Body_y[1785] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1786) begin
                        n_Body_x[1786] = c_Body_x[1785];
                        n_Body_y[1786] = c_Body_y[1785];
                    end else begin
                        n_Body_x[1786] = c_Body_x[c_Size-1];
                        n_Body_y[1786] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1787) begin
                        n_Body_x[1787] = c_Body_x[1786];
                        n_Body_y[1787] = c_Body_y[1786];
                    end else begin
                        n_Body_x[1787] = c_Body_x[c_Size-1];
                        n_Body_y[1787] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1788) begin
                        n_Body_x[1788] = c_Body_x[1787];
                        n_Body_y[1788] = c_Body_y[1787];
                    end else begin
                        n_Body_x[1788] = c_Body_x[c_Size-1];
                        n_Body_y[1788] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1789) begin
                        n_Body_x[1789] = c_Body_x[1788];
                        n_Body_y[1789] = c_Body_y[1788];
                    end else begin
                        n_Body_x[1789] = c_Body_x[c_Size-1];
                        n_Body_y[1789] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1790) begin
                        n_Body_x[1790] = c_Body_x[1789];
                        n_Body_y[1790] = c_Body_y[1789];
                    end else begin
                        n_Body_x[1790] = c_Body_x[c_Size-1];
                        n_Body_y[1790] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1791) begin
                        n_Body_x[1791] = c_Body_x[1790];
                        n_Body_y[1791] = c_Body_y[1790];
                    end else begin
                        n_Body_x[1791] = c_Body_x[c_Size-1];
                        n_Body_y[1791] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1792) begin
                        n_Body_x[1792] = c_Body_x[1791];
                        n_Body_y[1792] = c_Body_y[1791];
                    end else begin
                        n_Body_x[1792] = c_Body_x[c_Size-1];
                        n_Body_y[1792] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1793) begin
                        n_Body_x[1793] = c_Body_x[1792];
                        n_Body_y[1793] = c_Body_y[1792];
                    end else begin
                        n_Body_x[1793] = c_Body_x[c_Size-1];
                        n_Body_y[1793] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1794) begin
                        n_Body_x[1794] = c_Body_x[1793];
                        n_Body_y[1794] = c_Body_y[1793];
                    end else begin
                        n_Body_x[1794] = c_Body_x[c_Size-1];
                        n_Body_y[1794] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1795) begin
                        n_Body_x[1795] = c_Body_x[1794];
                        n_Body_y[1795] = c_Body_y[1794];
                    end else begin
                        n_Body_x[1795] = c_Body_x[c_Size-1];
                        n_Body_y[1795] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1796) begin
                        n_Body_x[1796] = c_Body_x[1795];
                        n_Body_y[1796] = c_Body_y[1795];
                    end else begin
                        n_Body_x[1796] = c_Body_x[c_Size-1];
                        n_Body_y[1796] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1797) begin
                        n_Body_x[1797] = c_Body_x[1796];
                        n_Body_y[1797] = c_Body_y[1796];
                    end else begin
                        n_Body_x[1797] = c_Body_x[c_Size-1];
                        n_Body_y[1797] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1798) begin
                        n_Body_x[1798] = c_Body_x[1797];
                        n_Body_y[1798] = c_Body_y[1797];
                    end else begin
                        n_Body_x[1798] = c_Body_x[c_Size-1];
                        n_Body_y[1798] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1799) begin
                        n_Body_x[1799] = c_Body_x[1798];
                        n_Body_y[1799] = c_Body_y[1798];
                    end else begin
                        n_Body_x[1799] = c_Body_x[c_Size-1];
                        n_Body_y[1799] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1800) begin
                        n_Body_x[1800] = c_Body_x[1799];
                        n_Body_y[1800] = c_Body_y[1799];
                    end else begin
                        n_Body_x[1800] = c_Body_x[c_Size-1];
                        n_Body_y[1800] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1801) begin
                        n_Body_x[1801] = c_Body_x[1800];
                        n_Body_y[1801] = c_Body_y[1800];
                    end else begin
                        n_Body_x[1801] = c_Body_x[c_Size-1];
                        n_Body_y[1801] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1802) begin
                        n_Body_x[1802] = c_Body_x[1801];
                        n_Body_y[1802] = c_Body_y[1801];
                    end else begin
                        n_Body_x[1802] = c_Body_x[c_Size-1];
                        n_Body_y[1802] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1803) begin
                        n_Body_x[1803] = c_Body_x[1802];
                        n_Body_y[1803] = c_Body_y[1802];
                    end else begin
                        n_Body_x[1803] = c_Body_x[c_Size-1];
                        n_Body_y[1803] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1804) begin
                        n_Body_x[1804] = c_Body_x[1803];
                        n_Body_y[1804] = c_Body_y[1803];
                    end else begin
                        n_Body_x[1804] = c_Body_x[c_Size-1];
                        n_Body_y[1804] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1805) begin
                        n_Body_x[1805] = c_Body_x[1804];
                        n_Body_y[1805] = c_Body_y[1804];
                    end else begin
                        n_Body_x[1805] = c_Body_x[c_Size-1];
                        n_Body_y[1805] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1806) begin
                        n_Body_x[1806] = c_Body_x[1805];
                        n_Body_y[1806] = c_Body_y[1805];
                    end else begin
                        n_Body_x[1806] = c_Body_x[c_Size-1];
                        n_Body_y[1806] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1807) begin
                        n_Body_x[1807] = c_Body_x[1806];
                        n_Body_y[1807] = c_Body_y[1806];
                    end else begin
                        n_Body_x[1807] = c_Body_x[c_Size-1];
                        n_Body_y[1807] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1808) begin
                        n_Body_x[1808] = c_Body_x[1807];
                        n_Body_y[1808] = c_Body_y[1807];
                    end else begin
                        n_Body_x[1808] = c_Body_x[c_Size-1];
                        n_Body_y[1808] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1809) begin
                        n_Body_x[1809] = c_Body_x[1808];
                        n_Body_y[1809] = c_Body_y[1808];
                    end else begin
                        n_Body_x[1809] = c_Body_x[c_Size-1];
                        n_Body_y[1809] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1810) begin
                        n_Body_x[1810] = c_Body_x[1809];
                        n_Body_y[1810] = c_Body_y[1809];
                    end else begin
                        n_Body_x[1810] = c_Body_x[c_Size-1];
                        n_Body_y[1810] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1811) begin
                        n_Body_x[1811] = c_Body_x[1810];
                        n_Body_y[1811] = c_Body_y[1810];
                    end else begin
                        n_Body_x[1811] = c_Body_x[c_Size-1];
                        n_Body_y[1811] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1812) begin
                        n_Body_x[1812] = c_Body_x[1811];
                        n_Body_y[1812] = c_Body_y[1811];
                    end else begin
                        n_Body_x[1812] = c_Body_x[c_Size-1];
                        n_Body_y[1812] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1813) begin
                        n_Body_x[1813] = c_Body_x[1812];
                        n_Body_y[1813] = c_Body_y[1812];
                    end else begin
                        n_Body_x[1813] = c_Body_x[c_Size-1];
                        n_Body_y[1813] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1814) begin
                        n_Body_x[1814] = c_Body_x[1813];
                        n_Body_y[1814] = c_Body_y[1813];
                    end else begin
                        n_Body_x[1814] = c_Body_x[c_Size-1];
                        n_Body_y[1814] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1815) begin
                        n_Body_x[1815] = c_Body_x[1814];
                        n_Body_y[1815] = c_Body_y[1814];
                    end else begin
                        n_Body_x[1815] = c_Body_x[c_Size-1];
                        n_Body_y[1815] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1816) begin
                        n_Body_x[1816] = c_Body_x[1815];
                        n_Body_y[1816] = c_Body_y[1815];
                    end else begin
                        n_Body_x[1816] = c_Body_x[c_Size-1];
                        n_Body_y[1816] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1817) begin
                        n_Body_x[1817] = c_Body_x[1816];
                        n_Body_y[1817] = c_Body_y[1816];
                    end else begin
                        n_Body_x[1817] = c_Body_x[c_Size-1];
                        n_Body_y[1817] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1818) begin
                        n_Body_x[1818] = c_Body_x[1817];
                        n_Body_y[1818] = c_Body_y[1817];
                    end else begin
                        n_Body_x[1818] = c_Body_x[c_Size-1];
                        n_Body_y[1818] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1819) begin
                        n_Body_x[1819] = c_Body_x[1818];
                        n_Body_y[1819] = c_Body_y[1818];
                    end else begin
                        n_Body_x[1819] = c_Body_x[c_Size-1];
                        n_Body_y[1819] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1820) begin
                        n_Body_x[1820] = c_Body_x[1819];
                        n_Body_y[1820] = c_Body_y[1819];
                    end else begin
                        n_Body_x[1820] = c_Body_x[c_Size-1];
                        n_Body_y[1820] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1821) begin
                        n_Body_x[1821] = c_Body_x[1820];
                        n_Body_y[1821] = c_Body_y[1820];
                    end else begin
                        n_Body_x[1821] = c_Body_x[c_Size-1];
                        n_Body_y[1821] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1822) begin
                        n_Body_x[1822] = c_Body_x[1821];
                        n_Body_y[1822] = c_Body_y[1821];
                    end else begin
                        n_Body_x[1822] = c_Body_x[c_Size-1];
                        n_Body_y[1822] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1823) begin
                        n_Body_x[1823] = c_Body_x[1822];
                        n_Body_y[1823] = c_Body_y[1822];
                    end else begin
                        n_Body_x[1823] = c_Body_x[c_Size-1];
                        n_Body_y[1823] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1824) begin
                        n_Body_x[1824] = c_Body_x[1823];
                        n_Body_y[1824] = c_Body_y[1823];
                    end else begin
                        n_Body_x[1824] = c_Body_x[c_Size-1];
                        n_Body_y[1824] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1825) begin
                        n_Body_x[1825] = c_Body_x[1824];
                        n_Body_y[1825] = c_Body_y[1824];
                    end else begin
                        n_Body_x[1825] = c_Body_x[c_Size-1];
                        n_Body_y[1825] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1826) begin
                        n_Body_x[1826] = c_Body_x[1825];
                        n_Body_y[1826] = c_Body_y[1825];
                    end else begin
                        n_Body_x[1826] = c_Body_x[c_Size-1];
                        n_Body_y[1826] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1827) begin
                        n_Body_x[1827] = c_Body_x[1826];
                        n_Body_y[1827] = c_Body_y[1826];
                    end else begin
                        n_Body_x[1827] = c_Body_x[c_Size-1];
                        n_Body_y[1827] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1828) begin
                        n_Body_x[1828] = c_Body_x[1827];
                        n_Body_y[1828] = c_Body_y[1827];
                    end else begin
                        n_Body_x[1828] = c_Body_x[c_Size-1];
                        n_Body_y[1828] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1829) begin
                        n_Body_x[1829] = c_Body_x[1828];
                        n_Body_y[1829] = c_Body_y[1828];
                    end else begin
                        n_Body_x[1829] = c_Body_x[c_Size-1];
                        n_Body_y[1829] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1830) begin
                        n_Body_x[1830] = c_Body_x[1829];
                        n_Body_y[1830] = c_Body_y[1829];
                    end else begin
                        n_Body_x[1830] = c_Body_x[c_Size-1];
                        n_Body_y[1830] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1831) begin
                        n_Body_x[1831] = c_Body_x[1830];
                        n_Body_y[1831] = c_Body_y[1830];
                    end else begin
                        n_Body_x[1831] = c_Body_x[c_Size-1];
                        n_Body_y[1831] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1832) begin
                        n_Body_x[1832] = c_Body_x[1831];
                        n_Body_y[1832] = c_Body_y[1831];
                    end else begin
                        n_Body_x[1832] = c_Body_x[c_Size-1];
                        n_Body_y[1832] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1833) begin
                        n_Body_x[1833] = c_Body_x[1832];
                        n_Body_y[1833] = c_Body_y[1832];
                    end else begin
                        n_Body_x[1833] = c_Body_x[c_Size-1];
                        n_Body_y[1833] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1834) begin
                        n_Body_x[1834] = c_Body_x[1833];
                        n_Body_y[1834] = c_Body_y[1833];
                    end else begin
                        n_Body_x[1834] = c_Body_x[c_Size-1];
                        n_Body_y[1834] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1835) begin
                        n_Body_x[1835] = c_Body_x[1834];
                        n_Body_y[1835] = c_Body_y[1834];
                    end else begin
                        n_Body_x[1835] = c_Body_x[c_Size-1];
                        n_Body_y[1835] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1836) begin
                        n_Body_x[1836] = c_Body_x[1835];
                        n_Body_y[1836] = c_Body_y[1835];
                    end else begin
                        n_Body_x[1836] = c_Body_x[c_Size-1];
                        n_Body_y[1836] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1837) begin
                        n_Body_x[1837] = c_Body_x[1836];
                        n_Body_y[1837] = c_Body_y[1836];
                    end else begin
                        n_Body_x[1837] = c_Body_x[c_Size-1];
                        n_Body_y[1837] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1838) begin
                        n_Body_x[1838] = c_Body_x[1837];
                        n_Body_y[1838] = c_Body_y[1837];
                    end else begin
                        n_Body_x[1838] = c_Body_x[c_Size-1];
                        n_Body_y[1838] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1839) begin
                        n_Body_x[1839] = c_Body_x[1838];
                        n_Body_y[1839] = c_Body_y[1838];
                    end else begin
                        n_Body_x[1839] = c_Body_x[c_Size-1];
                        n_Body_y[1839] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1840) begin
                        n_Body_x[1840] = c_Body_x[1839];
                        n_Body_y[1840] = c_Body_y[1839];
                    end else begin
                        n_Body_x[1840] = c_Body_x[c_Size-1];
                        n_Body_y[1840] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1841) begin
                        n_Body_x[1841] = c_Body_x[1840];
                        n_Body_y[1841] = c_Body_y[1840];
                    end else begin
                        n_Body_x[1841] = c_Body_x[c_Size-1];
                        n_Body_y[1841] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1842) begin
                        n_Body_x[1842] = c_Body_x[1841];
                        n_Body_y[1842] = c_Body_y[1841];
                    end else begin
                        n_Body_x[1842] = c_Body_x[c_Size-1];
                        n_Body_y[1842] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1843) begin
                        n_Body_x[1843] = c_Body_x[1842];
                        n_Body_y[1843] = c_Body_y[1842];
                    end else begin
                        n_Body_x[1843] = c_Body_x[c_Size-1];
                        n_Body_y[1843] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1844) begin
                        n_Body_x[1844] = c_Body_x[1843];
                        n_Body_y[1844] = c_Body_y[1843];
                    end else begin
                        n_Body_x[1844] = c_Body_x[c_Size-1];
                        n_Body_y[1844] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1845) begin
                        n_Body_x[1845] = c_Body_x[1844];
                        n_Body_y[1845] = c_Body_y[1844];
                    end else begin
                        n_Body_x[1845] = c_Body_x[c_Size-1];
                        n_Body_y[1845] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1846) begin
                        n_Body_x[1846] = c_Body_x[1845];
                        n_Body_y[1846] = c_Body_y[1845];
                    end else begin
                        n_Body_x[1846] = c_Body_x[c_Size-1];
                        n_Body_y[1846] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1847) begin
                        n_Body_x[1847] = c_Body_x[1846];
                        n_Body_y[1847] = c_Body_y[1846];
                    end else begin
                        n_Body_x[1847] = c_Body_x[c_Size-1];
                        n_Body_y[1847] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1848) begin
                        n_Body_x[1848] = c_Body_x[1847];
                        n_Body_y[1848] = c_Body_y[1847];
                    end else begin
                        n_Body_x[1848] = c_Body_x[c_Size-1];
                        n_Body_y[1848] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1849) begin
                        n_Body_x[1849] = c_Body_x[1848];
                        n_Body_y[1849] = c_Body_y[1848];
                    end else begin
                        n_Body_x[1849] = c_Body_x[c_Size-1];
                        n_Body_y[1849] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1850) begin
                        n_Body_x[1850] = c_Body_x[1849];
                        n_Body_y[1850] = c_Body_y[1849];
                    end else begin
                        n_Body_x[1850] = c_Body_x[c_Size-1];
                        n_Body_y[1850] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1851) begin
                        n_Body_x[1851] = c_Body_x[1850];
                        n_Body_y[1851] = c_Body_y[1850];
                    end else begin
                        n_Body_x[1851] = c_Body_x[c_Size-1];
                        n_Body_y[1851] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1852) begin
                        n_Body_x[1852] = c_Body_x[1851];
                        n_Body_y[1852] = c_Body_y[1851];
                    end else begin
                        n_Body_x[1852] = c_Body_x[c_Size-1];
                        n_Body_y[1852] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1853) begin
                        n_Body_x[1853] = c_Body_x[1852];
                        n_Body_y[1853] = c_Body_y[1852];
                    end else begin
                        n_Body_x[1853] = c_Body_x[c_Size-1];
                        n_Body_y[1853] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1854) begin
                        n_Body_x[1854] = c_Body_x[1853];
                        n_Body_y[1854] = c_Body_y[1853];
                    end else begin
                        n_Body_x[1854] = c_Body_x[c_Size-1];
                        n_Body_y[1854] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1855) begin
                        n_Body_x[1855] = c_Body_x[1854];
                        n_Body_y[1855] = c_Body_y[1854];
                    end else begin
                        n_Body_x[1855] = c_Body_x[c_Size-1];
                        n_Body_y[1855] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1856) begin
                        n_Body_x[1856] = c_Body_x[1855];
                        n_Body_y[1856] = c_Body_y[1855];
                    end else begin
                        n_Body_x[1856] = c_Body_x[c_Size-1];
                        n_Body_y[1856] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1857) begin
                        n_Body_x[1857] = c_Body_x[1856];
                        n_Body_y[1857] = c_Body_y[1856];
                    end else begin
                        n_Body_x[1857] = c_Body_x[c_Size-1];
                        n_Body_y[1857] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1858) begin
                        n_Body_x[1858] = c_Body_x[1857];
                        n_Body_y[1858] = c_Body_y[1857];
                    end else begin
                        n_Body_x[1858] = c_Body_x[c_Size-1];
                        n_Body_y[1858] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1859) begin
                        n_Body_x[1859] = c_Body_x[1858];
                        n_Body_y[1859] = c_Body_y[1858];
                    end else begin
                        n_Body_x[1859] = c_Body_x[c_Size-1];
                        n_Body_y[1859] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1860) begin
                        n_Body_x[1860] = c_Body_x[1859];
                        n_Body_y[1860] = c_Body_y[1859];
                    end else begin
                        n_Body_x[1860] = c_Body_x[c_Size-1];
                        n_Body_y[1860] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1861) begin
                        n_Body_x[1861] = c_Body_x[1860];
                        n_Body_y[1861] = c_Body_y[1860];
                    end else begin
                        n_Body_x[1861] = c_Body_x[c_Size-1];
                        n_Body_y[1861] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1862) begin
                        n_Body_x[1862] = c_Body_x[1861];
                        n_Body_y[1862] = c_Body_y[1861];
                    end else begin
                        n_Body_x[1862] = c_Body_x[c_Size-1];
                        n_Body_y[1862] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1863) begin
                        n_Body_x[1863] = c_Body_x[1862];
                        n_Body_y[1863] = c_Body_y[1862];
                    end else begin
                        n_Body_x[1863] = c_Body_x[c_Size-1];
                        n_Body_y[1863] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1864) begin
                        n_Body_x[1864] = c_Body_x[1863];
                        n_Body_y[1864] = c_Body_y[1863];
                    end else begin
                        n_Body_x[1864] = c_Body_x[c_Size-1];
                        n_Body_y[1864] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1865) begin
                        n_Body_x[1865] = c_Body_x[1864];
                        n_Body_y[1865] = c_Body_y[1864];
                    end else begin
                        n_Body_x[1865] = c_Body_x[c_Size-1];
                        n_Body_y[1865] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1866) begin
                        n_Body_x[1866] = c_Body_x[1865];
                        n_Body_y[1866] = c_Body_y[1865];
                    end else begin
                        n_Body_x[1866] = c_Body_x[c_Size-1];
                        n_Body_y[1866] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1867) begin
                        n_Body_x[1867] = c_Body_x[1866];
                        n_Body_y[1867] = c_Body_y[1866];
                    end else begin
                        n_Body_x[1867] = c_Body_x[c_Size-1];
                        n_Body_y[1867] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1868) begin
                        n_Body_x[1868] = c_Body_x[1867];
                        n_Body_y[1868] = c_Body_y[1867];
                    end else begin
                        n_Body_x[1868] = c_Body_x[c_Size-1];
                        n_Body_y[1868] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1869) begin
                        n_Body_x[1869] = c_Body_x[1868];
                        n_Body_y[1869] = c_Body_y[1868];
                    end else begin
                        n_Body_x[1869] = c_Body_x[c_Size-1];
                        n_Body_y[1869] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1870) begin
                        n_Body_x[1870] = c_Body_x[1869];
                        n_Body_y[1870] = c_Body_y[1869];
                    end else begin
                        n_Body_x[1870] = c_Body_x[c_Size-1];
                        n_Body_y[1870] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1871) begin
                        n_Body_x[1871] = c_Body_x[1870];
                        n_Body_y[1871] = c_Body_y[1870];
                    end else begin
                        n_Body_x[1871] = c_Body_x[c_Size-1];
                        n_Body_y[1871] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1872) begin
                        n_Body_x[1872] = c_Body_x[1871];
                        n_Body_y[1872] = c_Body_y[1871];
                    end else begin
                        n_Body_x[1872] = c_Body_x[c_Size-1];
                        n_Body_y[1872] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1873) begin
                        n_Body_x[1873] = c_Body_x[1872];
                        n_Body_y[1873] = c_Body_y[1872];
                    end else begin
                        n_Body_x[1873] = c_Body_x[c_Size-1];
                        n_Body_y[1873] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1874) begin
                        n_Body_x[1874] = c_Body_x[1873];
                        n_Body_y[1874] = c_Body_y[1873];
                    end else begin
                        n_Body_x[1874] = c_Body_x[c_Size-1];
                        n_Body_y[1874] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1875) begin
                        n_Body_x[1875] = c_Body_x[1874];
                        n_Body_y[1875] = c_Body_y[1874];
                    end else begin
                        n_Body_x[1875] = c_Body_x[c_Size-1];
                        n_Body_y[1875] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1876) begin
                        n_Body_x[1876] = c_Body_x[1875];
                        n_Body_y[1876] = c_Body_y[1875];
                    end else begin
                        n_Body_x[1876] = c_Body_x[c_Size-1];
                        n_Body_y[1876] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1877) begin
                        n_Body_x[1877] = c_Body_x[1876];
                        n_Body_y[1877] = c_Body_y[1876];
                    end else begin
                        n_Body_x[1877] = c_Body_x[c_Size-1];
                        n_Body_y[1877] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1878) begin
                        n_Body_x[1878] = c_Body_x[1877];
                        n_Body_y[1878] = c_Body_y[1877];
                    end else begin
                        n_Body_x[1878] = c_Body_x[c_Size-1];
                        n_Body_y[1878] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1879) begin
                        n_Body_x[1879] = c_Body_x[1878];
                        n_Body_y[1879] = c_Body_y[1878];
                    end else begin
                        n_Body_x[1879] = c_Body_x[c_Size-1];
                        n_Body_y[1879] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1880) begin
                        n_Body_x[1880] = c_Body_x[1879];
                        n_Body_y[1880] = c_Body_y[1879];
                    end else begin
                        n_Body_x[1880] = c_Body_x[c_Size-1];
                        n_Body_y[1880] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1881) begin
                        n_Body_x[1881] = c_Body_x[1880];
                        n_Body_y[1881] = c_Body_y[1880];
                    end else begin
                        n_Body_x[1881] = c_Body_x[c_Size-1];
                        n_Body_y[1881] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1882) begin
                        n_Body_x[1882] = c_Body_x[1881];
                        n_Body_y[1882] = c_Body_y[1881];
                    end else begin
                        n_Body_x[1882] = c_Body_x[c_Size-1];
                        n_Body_y[1882] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1883) begin
                        n_Body_x[1883] = c_Body_x[1882];
                        n_Body_y[1883] = c_Body_y[1882];
                    end else begin
                        n_Body_x[1883] = c_Body_x[c_Size-1];
                        n_Body_y[1883] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1884) begin
                        n_Body_x[1884] = c_Body_x[1883];
                        n_Body_y[1884] = c_Body_y[1883];
                    end else begin
                        n_Body_x[1884] = c_Body_x[c_Size-1];
                        n_Body_y[1884] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1885) begin
                        n_Body_x[1885] = c_Body_x[1884];
                        n_Body_y[1885] = c_Body_y[1884];
                    end else begin
                        n_Body_x[1885] = c_Body_x[c_Size-1];
                        n_Body_y[1885] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1886) begin
                        n_Body_x[1886] = c_Body_x[1885];
                        n_Body_y[1886] = c_Body_y[1885];
                    end else begin
                        n_Body_x[1886] = c_Body_x[c_Size-1];
                        n_Body_y[1886] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1887) begin
                        n_Body_x[1887] = c_Body_x[1886];
                        n_Body_y[1887] = c_Body_y[1886];
                    end else begin
                        n_Body_x[1887] = c_Body_x[c_Size-1];
                        n_Body_y[1887] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1888) begin
                        n_Body_x[1888] = c_Body_x[1887];
                        n_Body_y[1888] = c_Body_y[1887];
                    end else begin
                        n_Body_x[1888] = c_Body_x[c_Size-1];
                        n_Body_y[1888] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1889) begin
                        n_Body_x[1889] = c_Body_x[1888];
                        n_Body_y[1889] = c_Body_y[1888];
                    end else begin
                        n_Body_x[1889] = c_Body_x[c_Size-1];
                        n_Body_y[1889] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1890) begin
                        n_Body_x[1890] = c_Body_x[1889];
                        n_Body_y[1890] = c_Body_y[1889];
                    end else begin
                        n_Body_x[1890] = c_Body_x[c_Size-1];
                        n_Body_y[1890] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1891) begin
                        n_Body_x[1891] = c_Body_x[1890];
                        n_Body_y[1891] = c_Body_y[1890];
                    end else begin
                        n_Body_x[1891] = c_Body_x[c_Size-1];
                        n_Body_y[1891] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1892) begin
                        n_Body_x[1892] = c_Body_x[1891];
                        n_Body_y[1892] = c_Body_y[1891];
                    end else begin
                        n_Body_x[1892] = c_Body_x[c_Size-1];
                        n_Body_y[1892] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1893) begin
                        n_Body_x[1893] = c_Body_x[1892];
                        n_Body_y[1893] = c_Body_y[1892];
                    end else begin
                        n_Body_x[1893] = c_Body_x[c_Size-1];
                        n_Body_y[1893] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1894) begin
                        n_Body_x[1894] = c_Body_x[1893];
                        n_Body_y[1894] = c_Body_y[1893];
                    end else begin
                        n_Body_x[1894] = c_Body_x[c_Size-1];
                        n_Body_y[1894] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1895) begin
                        n_Body_x[1895] = c_Body_x[1894];
                        n_Body_y[1895] = c_Body_y[1894];
                    end else begin
                        n_Body_x[1895] = c_Body_x[c_Size-1];
                        n_Body_y[1895] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1896) begin
                        n_Body_x[1896] = c_Body_x[1895];
                        n_Body_y[1896] = c_Body_y[1895];
                    end else begin
                        n_Body_x[1896] = c_Body_x[c_Size-1];
                        n_Body_y[1896] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1897) begin
                        n_Body_x[1897] = c_Body_x[1896];
                        n_Body_y[1897] = c_Body_y[1896];
                    end else begin
                        n_Body_x[1897] = c_Body_x[c_Size-1];
                        n_Body_y[1897] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1898) begin
                        n_Body_x[1898] = c_Body_x[1897];
                        n_Body_y[1898] = c_Body_y[1897];
                    end else begin
                        n_Body_x[1898] = c_Body_x[c_Size-1];
                        n_Body_y[1898] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1899) begin
                        n_Body_x[1899] = c_Body_x[1898];
                        n_Body_y[1899] = c_Body_y[1898];
                    end else begin
                        n_Body_x[1899] = c_Body_x[c_Size-1];
                        n_Body_y[1899] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1900) begin
                        n_Body_x[1900] = c_Body_x[1899];
                        n_Body_y[1900] = c_Body_y[1899];
                    end else begin
                        n_Body_x[1900] = c_Body_x[c_Size-1];
                        n_Body_y[1900] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1901) begin
                        n_Body_x[1901] = c_Body_x[1900];
                        n_Body_y[1901] = c_Body_y[1900];
                    end else begin
                        n_Body_x[1901] = c_Body_x[c_Size-1];
                        n_Body_y[1901] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1902) begin
                        n_Body_x[1902] = c_Body_x[1901];
                        n_Body_y[1902] = c_Body_y[1901];
                    end else begin
                        n_Body_x[1902] = c_Body_x[c_Size-1];
                        n_Body_y[1902] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1903) begin
                        n_Body_x[1903] = c_Body_x[1902];
                        n_Body_y[1903] = c_Body_y[1902];
                    end else begin
                        n_Body_x[1903] = c_Body_x[c_Size-1];
                        n_Body_y[1903] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1904) begin
                        n_Body_x[1904] = c_Body_x[1903];
                        n_Body_y[1904] = c_Body_y[1903];
                    end else begin
                        n_Body_x[1904] = c_Body_x[c_Size-1];
                        n_Body_y[1904] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1905) begin
                        n_Body_x[1905] = c_Body_x[1904];
                        n_Body_y[1905] = c_Body_y[1904];
                    end else begin
                        n_Body_x[1905] = c_Body_x[c_Size-1];
                        n_Body_y[1905] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1906) begin
                        n_Body_x[1906] = c_Body_x[1905];
                        n_Body_y[1906] = c_Body_y[1905];
                    end else begin
                        n_Body_x[1906] = c_Body_x[c_Size-1];
                        n_Body_y[1906] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1907) begin
                        n_Body_x[1907] = c_Body_x[1906];
                        n_Body_y[1907] = c_Body_y[1906];
                    end else begin
                        n_Body_x[1907] = c_Body_x[c_Size-1];
                        n_Body_y[1907] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1908) begin
                        n_Body_x[1908] = c_Body_x[1907];
                        n_Body_y[1908] = c_Body_y[1907];
                    end else begin
                        n_Body_x[1908] = c_Body_x[c_Size-1];
                        n_Body_y[1908] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1909) begin
                        n_Body_x[1909] = c_Body_x[1908];
                        n_Body_y[1909] = c_Body_y[1908];
                    end else begin
                        n_Body_x[1909] = c_Body_x[c_Size-1];
                        n_Body_y[1909] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1910) begin
                        n_Body_x[1910] = c_Body_x[1909];
                        n_Body_y[1910] = c_Body_y[1909];
                    end else begin
                        n_Body_x[1910] = c_Body_x[c_Size-1];
                        n_Body_y[1910] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1911) begin
                        n_Body_x[1911] = c_Body_x[1910];
                        n_Body_y[1911] = c_Body_y[1910];
                    end else begin
                        n_Body_x[1911] = c_Body_x[c_Size-1];
                        n_Body_y[1911] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1912) begin
                        n_Body_x[1912] = c_Body_x[1911];
                        n_Body_y[1912] = c_Body_y[1911];
                    end else begin
                        n_Body_x[1912] = c_Body_x[c_Size-1];
                        n_Body_y[1912] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1913) begin
                        n_Body_x[1913] = c_Body_x[1912];
                        n_Body_y[1913] = c_Body_y[1912];
                    end else begin
                        n_Body_x[1913] = c_Body_x[c_Size-1];
                        n_Body_y[1913] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1914) begin
                        n_Body_x[1914] = c_Body_x[1913];
                        n_Body_y[1914] = c_Body_y[1913];
                    end else begin
                        n_Body_x[1914] = c_Body_x[c_Size-1];
                        n_Body_y[1914] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1915) begin
                        n_Body_x[1915] = c_Body_x[1914];
                        n_Body_y[1915] = c_Body_y[1914];
                    end else begin
                        n_Body_x[1915] = c_Body_x[c_Size-1];
                        n_Body_y[1915] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1916) begin
                        n_Body_x[1916] = c_Body_x[1915];
                        n_Body_y[1916] = c_Body_y[1915];
                    end else begin
                        n_Body_x[1916] = c_Body_x[c_Size-1];
                        n_Body_y[1916] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1917) begin
                        n_Body_x[1917] = c_Body_x[1916];
                        n_Body_y[1917] = c_Body_y[1916];
                    end else begin
                        n_Body_x[1917] = c_Body_x[c_Size-1];
                        n_Body_y[1917] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1918) begin
                        n_Body_x[1918] = c_Body_x[1917];
                        n_Body_y[1918] = c_Body_y[1917];
                    end else begin
                        n_Body_x[1918] = c_Body_x[c_Size-1];
                        n_Body_y[1918] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1919) begin
                        n_Body_x[1919] = c_Body_x[1918];
                        n_Body_y[1919] = c_Body_y[1918];
                    end else begin
                        n_Body_x[1919] = c_Body_x[c_Size-1];
                        n_Body_y[1919] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1920) begin
                        n_Body_x[1920] = c_Body_x[1919];
                        n_Body_y[1920] = c_Body_y[1919];
                    end else begin
                        n_Body_x[1920] = c_Body_x[c_Size-1];
                        n_Body_y[1920] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1921) begin
                        n_Body_x[1921] = c_Body_x[1920];
                        n_Body_y[1921] = c_Body_y[1920];
                    end else begin
                        n_Body_x[1921] = c_Body_x[c_Size-1];
                        n_Body_y[1921] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1922) begin
                        n_Body_x[1922] = c_Body_x[1921];
                        n_Body_y[1922] = c_Body_y[1921];
                    end else begin
                        n_Body_x[1922] = c_Body_x[c_Size-1];
                        n_Body_y[1922] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1923) begin
                        n_Body_x[1923] = c_Body_x[1922];
                        n_Body_y[1923] = c_Body_y[1922];
                    end else begin
                        n_Body_x[1923] = c_Body_x[c_Size-1];
                        n_Body_y[1923] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1924) begin
                        n_Body_x[1924] = c_Body_x[1923];
                        n_Body_y[1924] = c_Body_y[1923];
                    end else begin
                        n_Body_x[1924] = c_Body_x[c_Size-1];
                        n_Body_y[1924] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1925) begin
                        n_Body_x[1925] = c_Body_x[1924];
                        n_Body_y[1925] = c_Body_y[1924];
                    end else begin
                        n_Body_x[1925] = c_Body_x[c_Size-1];
                        n_Body_y[1925] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1926) begin
                        n_Body_x[1926] = c_Body_x[1925];
                        n_Body_y[1926] = c_Body_y[1925];
                    end else begin
                        n_Body_x[1926] = c_Body_x[c_Size-1];
                        n_Body_y[1926] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1927) begin
                        n_Body_x[1927] = c_Body_x[1926];
                        n_Body_y[1927] = c_Body_y[1926];
                    end else begin
                        n_Body_x[1927] = c_Body_x[c_Size-1];
                        n_Body_y[1927] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1928) begin
                        n_Body_x[1928] = c_Body_x[1927];
                        n_Body_y[1928] = c_Body_y[1927];
                    end else begin
                        n_Body_x[1928] = c_Body_x[c_Size-1];
                        n_Body_y[1928] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1929) begin
                        n_Body_x[1929] = c_Body_x[1928];
                        n_Body_y[1929] = c_Body_y[1928];
                    end else begin
                        n_Body_x[1929] = c_Body_x[c_Size-1];
                        n_Body_y[1929] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1930) begin
                        n_Body_x[1930] = c_Body_x[1929];
                        n_Body_y[1930] = c_Body_y[1929];
                    end else begin
                        n_Body_x[1930] = c_Body_x[c_Size-1];
                        n_Body_y[1930] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1931) begin
                        n_Body_x[1931] = c_Body_x[1930];
                        n_Body_y[1931] = c_Body_y[1930];
                    end else begin
                        n_Body_x[1931] = c_Body_x[c_Size-1];
                        n_Body_y[1931] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1932) begin
                        n_Body_x[1932] = c_Body_x[1931];
                        n_Body_y[1932] = c_Body_y[1931];
                    end else begin
                        n_Body_x[1932] = c_Body_x[c_Size-1];
                        n_Body_y[1932] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1933) begin
                        n_Body_x[1933] = c_Body_x[1932];
                        n_Body_y[1933] = c_Body_y[1932];
                    end else begin
                        n_Body_x[1933] = c_Body_x[c_Size-1];
                        n_Body_y[1933] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1934) begin
                        n_Body_x[1934] = c_Body_x[1933];
                        n_Body_y[1934] = c_Body_y[1933];
                    end else begin
                        n_Body_x[1934] = c_Body_x[c_Size-1];
                        n_Body_y[1934] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1935) begin
                        n_Body_x[1935] = c_Body_x[1934];
                        n_Body_y[1935] = c_Body_y[1934];
                    end else begin
                        n_Body_x[1935] = c_Body_x[c_Size-1];
                        n_Body_y[1935] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1936) begin
                        n_Body_x[1936] = c_Body_x[1935];
                        n_Body_y[1936] = c_Body_y[1935];
                    end else begin
                        n_Body_x[1936] = c_Body_x[c_Size-1];
                        n_Body_y[1936] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1937) begin
                        n_Body_x[1937] = c_Body_x[1936];
                        n_Body_y[1937] = c_Body_y[1936];
                    end else begin
                        n_Body_x[1937] = c_Body_x[c_Size-1];
                        n_Body_y[1937] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1938) begin
                        n_Body_x[1938] = c_Body_x[1937];
                        n_Body_y[1938] = c_Body_y[1937];
                    end else begin
                        n_Body_x[1938] = c_Body_x[c_Size-1];
                        n_Body_y[1938] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1939) begin
                        n_Body_x[1939] = c_Body_x[1938];
                        n_Body_y[1939] = c_Body_y[1938];
                    end else begin
                        n_Body_x[1939] = c_Body_x[c_Size-1];
                        n_Body_y[1939] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1940) begin
                        n_Body_x[1940] = c_Body_x[1939];
                        n_Body_y[1940] = c_Body_y[1939];
                    end else begin
                        n_Body_x[1940] = c_Body_x[c_Size-1];
                        n_Body_y[1940] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1941) begin
                        n_Body_x[1941] = c_Body_x[1940];
                        n_Body_y[1941] = c_Body_y[1940];
                    end else begin
                        n_Body_x[1941] = c_Body_x[c_Size-1];
                        n_Body_y[1941] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1942) begin
                        n_Body_x[1942] = c_Body_x[1941];
                        n_Body_y[1942] = c_Body_y[1941];
                    end else begin
                        n_Body_x[1942] = c_Body_x[c_Size-1];
                        n_Body_y[1942] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1943) begin
                        n_Body_x[1943] = c_Body_x[1942];
                        n_Body_y[1943] = c_Body_y[1942];
                    end else begin
                        n_Body_x[1943] = c_Body_x[c_Size-1];
                        n_Body_y[1943] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1944) begin
                        n_Body_x[1944] = c_Body_x[1943];
                        n_Body_y[1944] = c_Body_y[1943];
                    end else begin
                        n_Body_x[1944] = c_Body_x[c_Size-1];
                        n_Body_y[1944] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1945) begin
                        n_Body_x[1945] = c_Body_x[1944];
                        n_Body_y[1945] = c_Body_y[1944];
                    end else begin
                        n_Body_x[1945] = c_Body_x[c_Size-1];
                        n_Body_y[1945] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1946) begin
                        n_Body_x[1946] = c_Body_x[1945];
                        n_Body_y[1946] = c_Body_y[1945];
                    end else begin
                        n_Body_x[1946] = c_Body_x[c_Size-1];
                        n_Body_y[1946] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1947) begin
                        n_Body_x[1947] = c_Body_x[1946];
                        n_Body_y[1947] = c_Body_y[1946];
                    end else begin
                        n_Body_x[1947] = c_Body_x[c_Size-1];
                        n_Body_y[1947] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1948) begin
                        n_Body_x[1948] = c_Body_x[1947];
                        n_Body_y[1948] = c_Body_y[1947];
                    end else begin
                        n_Body_x[1948] = c_Body_x[c_Size-1];
                        n_Body_y[1948] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1949) begin
                        n_Body_x[1949] = c_Body_x[1948];
                        n_Body_y[1949] = c_Body_y[1948];
                    end else begin
                        n_Body_x[1949] = c_Body_x[c_Size-1];
                        n_Body_y[1949] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1950) begin
                        n_Body_x[1950] = c_Body_x[1949];
                        n_Body_y[1950] = c_Body_y[1949];
                    end else begin
                        n_Body_x[1950] = c_Body_x[c_Size-1];
                        n_Body_y[1950] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1951) begin
                        n_Body_x[1951] = c_Body_x[1950];
                        n_Body_y[1951] = c_Body_y[1950];
                    end else begin
                        n_Body_x[1951] = c_Body_x[c_Size-1];
                        n_Body_y[1951] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1952) begin
                        n_Body_x[1952] = c_Body_x[1951];
                        n_Body_y[1952] = c_Body_y[1951];
                    end else begin
                        n_Body_x[1952] = c_Body_x[c_Size-1];
                        n_Body_y[1952] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1953) begin
                        n_Body_x[1953] = c_Body_x[1952];
                        n_Body_y[1953] = c_Body_y[1952];
                    end else begin
                        n_Body_x[1953] = c_Body_x[c_Size-1];
                        n_Body_y[1953] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1954) begin
                        n_Body_x[1954] = c_Body_x[1953];
                        n_Body_y[1954] = c_Body_y[1953];
                    end else begin
                        n_Body_x[1954] = c_Body_x[c_Size-1];
                        n_Body_y[1954] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1955) begin
                        n_Body_x[1955] = c_Body_x[1954];
                        n_Body_y[1955] = c_Body_y[1954];
                    end else begin
                        n_Body_x[1955] = c_Body_x[c_Size-1];
                        n_Body_y[1955] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1956) begin
                        n_Body_x[1956] = c_Body_x[1955];
                        n_Body_y[1956] = c_Body_y[1955];
                    end else begin
                        n_Body_x[1956] = c_Body_x[c_Size-1];
                        n_Body_y[1956] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1957) begin
                        n_Body_x[1957] = c_Body_x[1956];
                        n_Body_y[1957] = c_Body_y[1956];
                    end else begin
                        n_Body_x[1957] = c_Body_x[c_Size-1];
                        n_Body_y[1957] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1958) begin
                        n_Body_x[1958] = c_Body_x[1957];
                        n_Body_y[1958] = c_Body_y[1957];
                    end else begin
                        n_Body_x[1958] = c_Body_x[c_Size-1];
                        n_Body_y[1958] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1959) begin
                        n_Body_x[1959] = c_Body_x[1958];
                        n_Body_y[1959] = c_Body_y[1958];
                    end else begin
                        n_Body_x[1959] = c_Body_x[c_Size-1];
                        n_Body_y[1959] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1960) begin
                        n_Body_x[1960] = c_Body_x[1959];
                        n_Body_y[1960] = c_Body_y[1959];
                    end else begin
                        n_Body_x[1960] = c_Body_x[c_Size-1];
                        n_Body_y[1960] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1961) begin
                        n_Body_x[1961] = c_Body_x[1960];
                        n_Body_y[1961] = c_Body_y[1960];
                    end else begin
                        n_Body_x[1961] = c_Body_x[c_Size-1];
                        n_Body_y[1961] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1962) begin
                        n_Body_x[1962] = c_Body_x[1961];
                        n_Body_y[1962] = c_Body_y[1961];
                    end else begin
                        n_Body_x[1962] = c_Body_x[c_Size-1];
                        n_Body_y[1962] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1963) begin
                        n_Body_x[1963] = c_Body_x[1962];
                        n_Body_y[1963] = c_Body_y[1962];
                    end else begin
                        n_Body_x[1963] = c_Body_x[c_Size-1];
                        n_Body_y[1963] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1964) begin
                        n_Body_x[1964] = c_Body_x[1963];
                        n_Body_y[1964] = c_Body_y[1963];
                    end else begin
                        n_Body_x[1964] = c_Body_x[c_Size-1];
                        n_Body_y[1964] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1965) begin
                        n_Body_x[1965] = c_Body_x[1964];
                        n_Body_y[1965] = c_Body_y[1964];
                    end else begin
                        n_Body_x[1965] = c_Body_x[c_Size-1];
                        n_Body_y[1965] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1966) begin
                        n_Body_x[1966] = c_Body_x[1965];
                        n_Body_y[1966] = c_Body_y[1965];
                    end else begin
                        n_Body_x[1966] = c_Body_x[c_Size-1];
                        n_Body_y[1966] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1967) begin
                        n_Body_x[1967] = c_Body_x[1966];
                        n_Body_y[1967] = c_Body_y[1966];
                    end else begin
                        n_Body_x[1967] = c_Body_x[c_Size-1];
                        n_Body_y[1967] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1968) begin
                        n_Body_x[1968] = c_Body_x[1967];
                        n_Body_y[1968] = c_Body_y[1967];
                    end else begin
                        n_Body_x[1968] = c_Body_x[c_Size-1];
                        n_Body_y[1968] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1969) begin
                        n_Body_x[1969] = c_Body_x[1968];
                        n_Body_y[1969] = c_Body_y[1968];
                    end else begin
                        n_Body_x[1969] = c_Body_x[c_Size-1];
                        n_Body_y[1969] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1970) begin
                        n_Body_x[1970] = c_Body_x[1969];
                        n_Body_y[1970] = c_Body_y[1969];
                    end else begin
                        n_Body_x[1970] = c_Body_x[c_Size-1];
                        n_Body_y[1970] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1971) begin
                        n_Body_x[1971] = c_Body_x[1970];
                        n_Body_y[1971] = c_Body_y[1970];
                    end else begin
                        n_Body_x[1971] = c_Body_x[c_Size-1];
                        n_Body_y[1971] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1972) begin
                        n_Body_x[1972] = c_Body_x[1971];
                        n_Body_y[1972] = c_Body_y[1971];
                    end else begin
                        n_Body_x[1972] = c_Body_x[c_Size-1];
                        n_Body_y[1972] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1973) begin
                        n_Body_x[1973] = c_Body_x[1972];
                        n_Body_y[1973] = c_Body_y[1972];
                    end else begin
                        n_Body_x[1973] = c_Body_x[c_Size-1];
                        n_Body_y[1973] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1974) begin
                        n_Body_x[1974] = c_Body_x[1973];
                        n_Body_y[1974] = c_Body_y[1973];
                    end else begin
                        n_Body_x[1974] = c_Body_x[c_Size-1];
                        n_Body_y[1974] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1975) begin
                        n_Body_x[1975] = c_Body_x[1974];
                        n_Body_y[1975] = c_Body_y[1974];
                    end else begin
                        n_Body_x[1975] = c_Body_x[c_Size-1];
                        n_Body_y[1975] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1976) begin
                        n_Body_x[1976] = c_Body_x[1975];
                        n_Body_y[1976] = c_Body_y[1975];
                    end else begin
                        n_Body_x[1976] = c_Body_x[c_Size-1];
                        n_Body_y[1976] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1977) begin
                        n_Body_x[1977] = c_Body_x[1976];
                        n_Body_y[1977] = c_Body_y[1976];
                    end else begin
                        n_Body_x[1977] = c_Body_x[c_Size-1];
                        n_Body_y[1977] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1978) begin
                        n_Body_x[1978] = c_Body_x[1977];
                        n_Body_y[1978] = c_Body_y[1977];
                    end else begin
                        n_Body_x[1978] = c_Body_x[c_Size-1];
                        n_Body_y[1978] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1979) begin
                        n_Body_x[1979] = c_Body_x[1978];
                        n_Body_y[1979] = c_Body_y[1978];
                    end else begin
                        n_Body_x[1979] = c_Body_x[c_Size-1];
                        n_Body_y[1979] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1980) begin
                        n_Body_x[1980] = c_Body_x[1979];
                        n_Body_y[1980] = c_Body_y[1979];
                    end else begin
                        n_Body_x[1980] = c_Body_x[c_Size-1];
                        n_Body_y[1980] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1981) begin
                        n_Body_x[1981] = c_Body_x[1980];
                        n_Body_y[1981] = c_Body_y[1980];
                    end else begin
                        n_Body_x[1981] = c_Body_x[c_Size-1];
                        n_Body_y[1981] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1982) begin
                        n_Body_x[1982] = c_Body_x[1981];
                        n_Body_y[1982] = c_Body_y[1981];
                    end else begin
                        n_Body_x[1982] = c_Body_x[c_Size-1];
                        n_Body_y[1982] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1983) begin
                        n_Body_x[1983] = c_Body_x[1982];
                        n_Body_y[1983] = c_Body_y[1982];
                    end else begin
                        n_Body_x[1983] = c_Body_x[c_Size-1];
                        n_Body_y[1983] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1984) begin
                        n_Body_x[1984] = c_Body_x[1983];
                        n_Body_y[1984] = c_Body_y[1983];
                    end else begin
                        n_Body_x[1984] = c_Body_x[c_Size-1];
                        n_Body_y[1984] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1985) begin
                        n_Body_x[1985] = c_Body_x[1984];
                        n_Body_y[1985] = c_Body_y[1984];
                    end else begin
                        n_Body_x[1985] = c_Body_x[c_Size-1];
                        n_Body_y[1985] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1986) begin
                        n_Body_x[1986] = c_Body_x[1985];
                        n_Body_y[1986] = c_Body_y[1985];
                    end else begin
                        n_Body_x[1986] = c_Body_x[c_Size-1];
                        n_Body_y[1986] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1987) begin
                        n_Body_x[1987] = c_Body_x[1986];
                        n_Body_y[1987] = c_Body_y[1986];
                    end else begin
                        n_Body_x[1987] = c_Body_x[c_Size-1];
                        n_Body_y[1987] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1988) begin
                        n_Body_x[1988] = c_Body_x[1987];
                        n_Body_y[1988] = c_Body_y[1987];
                    end else begin
                        n_Body_x[1988] = c_Body_x[c_Size-1];
                        n_Body_y[1988] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1989) begin
                        n_Body_x[1989] = c_Body_x[1988];
                        n_Body_y[1989] = c_Body_y[1988];
                    end else begin
                        n_Body_x[1989] = c_Body_x[c_Size-1];
                        n_Body_y[1989] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1990) begin
                        n_Body_x[1990] = c_Body_x[1989];
                        n_Body_y[1990] = c_Body_y[1989];
                    end else begin
                        n_Body_x[1990] = c_Body_x[c_Size-1];
                        n_Body_y[1990] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1991) begin
                        n_Body_x[1991] = c_Body_x[1990];
                        n_Body_y[1991] = c_Body_y[1990];
                    end else begin
                        n_Body_x[1991] = c_Body_x[c_Size-1];
                        n_Body_y[1991] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1992) begin
                        n_Body_x[1992] = c_Body_x[1991];
                        n_Body_y[1992] = c_Body_y[1991];
                    end else begin
                        n_Body_x[1992] = c_Body_x[c_Size-1];
                        n_Body_y[1992] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1993) begin
                        n_Body_x[1993] = c_Body_x[1992];
                        n_Body_y[1993] = c_Body_y[1992];
                    end else begin
                        n_Body_x[1993] = c_Body_x[c_Size-1];
                        n_Body_y[1993] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1994) begin
                        n_Body_x[1994] = c_Body_x[1993];
                        n_Body_y[1994] = c_Body_y[1993];
                    end else begin
                        n_Body_x[1994] = c_Body_x[c_Size-1];
                        n_Body_y[1994] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1995) begin
                        n_Body_x[1995] = c_Body_x[1994];
                        n_Body_y[1995] = c_Body_y[1994];
                    end else begin
                        n_Body_x[1995] = c_Body_x[c_Size-1];
                        n_Body_y[1995] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1996) begin
                        n_Body_x[1996] = c_Body_x[1995];
                        n_Body_y[1996] = c_Body_y[1995];
                    end else begin
                        n_Body_x[1996] = c_Body_x[c_Size-1];
                        n_Body_y[1996] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1997) begin
                        n_Body_x[1997] = c_Body_x[1996];
                        n_Body_y[1997] = c_Body_y[1996];
                    end else begin
                        n_Body_x[1997] = c_Body_x[c_Size-1];
                        n_Body_y[1997] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1998) begin
                        n_Body_x[1998] = c_Body_x[1997];
                        n_Body_y[1998] = c_Body_y[1997];
                    end else begin
                        n_Body_x[1998] = c_Body_x[c_Size-1];
                        n_Body_y[1998] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 1999) begin
                        n_Body_x[1999] = c_Body_x[1998];
                        n_Body_y[1999] = c_Body_y[1998];
                    end else begin
                        n_Body_x[1999] = c_Body_x[c_Size-1];
                        n_Body_y[1999] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2000) begin
                        n_Body_x[2000] = c_Body_x[1999];
                        n_Body_y[2000] = c_Body_y[1999];
                    end else begin
                        n_Body_x[2000] = c_Body_x[c_Size-1];
                        n_Body_y[2000] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2001) begin
                        n_Body_x[2001] = c_Body_x[2000];
                        n_Body_y[2001] = c_Body_y[2000];
                    end else begin
                        n_Body_x[2001] = c_Body_x[c_Size-1];
                        n_Body_y[2001] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2002) begin
                        n_Body_x[2002] = c_Body_x[2001];
                        n_Body_y[2002] = c_Body_y[2001];
                    end else begin
                        n_Body_x[2002] = c_Body_x[c_Size-1];
                        n_Body_y[2002] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2003) begin
                        n_Body_x[2003] = c_Body_x[2002];
                        n_Body_y[2003] = c_Body_y[2002];
                    end else begin
                        n_Body_x[2003] = c_Body_x[c_Size-1];
                        n_Body_y[2003] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2004) begin
                        n_Body_x[2004] = c_Body_x[2003];
                        n_Body_y[2004] = c_Body_y[2003];
                    end else begin
                        n_Body_x[2004] = c_Body_x[c_Size-1];
                        n_Body_y[2004] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2005) begin
                        n_Body_x[2005] = c_Body_x[2004];
                        n_Body_y[2005] = c_Body_y[2004];
                    end else begin
                        n_Body_x[2005] = c_Body_x[c_Size-1];
                        n_Body_y[2005] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2006) begin
                        n_Body_x[2006] = c_Body_x[2005];
                        n_Body_y[2006] = c_Body_y[2005];
                    end else begin
                        n_Body_x[2006] = c_Body_x[c_Size-1];
                        n_Body_y[2006] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2007) begin
                        n_Body_x[2007] = c_Body_x[2006];
                        n_Body_y[2007] = c_Body_y[2006];
                    end else begin
                        n_Body_x[2007] = c_Body_x[c_Size-1];
                        n_Body_y[2007] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2008) begin
                        n_Body_x[2008] = c_Body_x[2007];
                        n_Body_y[2008] = c_Body_y[2007];
                    end else begin
                        n_Body_x[2008] = c_Body_x[c_Size-1];
                        n_Body_y[2008] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2009) begin
                        n_Body_x[2009] = c_Body_x[2008];
                        n_Body_y[2009] = c_Body_y[2008];
                    end else begin
                        n_Body_x[2009] = c_Body_x[c_Size-1];
                        n_Body_y[2009] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2010) begin
                        n_Body_x[2010] = c_Body_x[2009];
                        n_Body_y[2010] = c_Body_y[2009];
                    end else begin
                        n_Body_x[2010] = c_Body_x[c_Size-1];
                        n_Body_y[2010] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2011) begin
                        n_Body_x[2011] = c_Body_x[2010];
                        n_Body_y[2011] = c_Body_y[2010];
                    end else begin
                        n_Body_x[2011] = c_Body_x[c_Size-1];
                        n_Body_y[2011] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2012) begin
                        n_Body_x[2012] = c_Body_x[2011];
                        n_Body_y[2012] = c_Body_y[2011];
                    end else begin
                        n_Body_x[2012] = c_Body_x[c_Size-1];
                        n_Body_y[2012] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2013) begin
                        n_Body_x[2013] = c_Body_x[2012];
                        n_Body_y[2013] = c_Body_y[2012];
                    end else begin
                        n_Body_x[2013] = c_Body_x[c_Size-1];
                        n_Body_y[2013] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2014) begin
                        n_Body_x[2014] = c_Body_x[2013];
                        n_Body_y[2014] = c_Body_y[2013];
                    end else begin
                        n_Body_x[2014] = c_Body_x[c_Size-1];
                        n_Body_y[2014] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2015) begin
                        n_Body_x[2015] = c_Body_x[2014];
                        n_Body_y[2015] = c_Body_y[2014];
                    end else begin
                        n_Body_x[2015] = c_Body_x[c_Size-1];
                        n_Body_y[2015] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2016) begin
                        n_Body_x[2016] = c_Body_x[2015];
                        n_Body_y[2016] = c_Body_y[2015];
                    end else begin
                        n_Body_x[2016] = c_Body_x[c_Size-1];
                        n_Body_y[2016] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2017) begin
                        n_Body_x[2017] = c_Body_x[2016];
                        n_Body_y[2017] = c_Body_y[2016];
                    end else begin
                        n_Body_x[2017] = c_Body_x[c_Size-1];
                        n_Body_y[2017] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2018) begin
                        n_Body_x[2018] = c_Body_x[2017];
                        n_Body_y[2018] = c_Body_y[2017];
                    end else begin
                        n_Body_x[2018] = c_Body_x[c_Size-1];
                        n_Body_y[2018] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2019) begin
                        n_Body_x[2019] = c_Body_x[2018];
                        n_Body_y[2019] = c_Body_y[2018];
                    end else begin
                        n_Body_x[2019] = c_Body_x[c_Size-1];
                        n_Body_y[2019] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2020) begin
                        n_Body_x[2020] = c_Body_x[2019];
                        n_Body_y[2020] = c_Body_y[2019];
                    end else begin
                        n_Body_x[2020] = c_Body_x[c_Size-1];
                        n_Body_y[2020] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2021) begin
                        n_Body_x[2021] = c_Body_x[2020];
                        n_Body_y[2021] = c_Body_y[2020];
                    end else begin
                        n_Body_x[2021] = c_Body_x[c_Size-1];
                        n_Body_y[2021] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2022) begin
                        n_Body_x[2022] = c_Body_x[2021];
                        n_Body_y[2022] = c_Body_y[2021];
                    end else begin
                        n_Body_x[2022] = c_Body_x[c_Size-1];
                        n_Body_y[2022] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2023) begin
                        n_Body_x[2023] = c_Body_x[2022];
                        n_Body_y[2023] = c_Body_y[2022];
                    end else begin
                        n_Body_x[2023] = c_Body_x[c_Size-1];
                        n_Body_y[2023] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2024) begin
                        n_Body_x[2024] = c_Body_x[2023];
                        n_Body_y[2024] = c_Body_y[2023];
                    end else begin
                        n_Body_x[2024] = c_Body_x[c_Size-1];
                        n_Body_y[2024] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2025) begin
                        n_Body_x[2025] = c_Body_x[2024];
                        n_Body_y[2025] = c_Body_y[2024];
                    end else begin
                        n_Body_x[2025] = c_Body_x[c_Size-1];
                        n_Body_y[2025] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2026) begin
                        n_Body_x[2026] = c_Body_x[2025];
                        n_Body_y[2026] = c_Body_y[2025];
                    end else begin
                        n_Body_x[2026] = c_Body_x[c_Size-1];
                        n_Body_y[2026] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2027) begin
                        n_Body_x[2027] = c_Body_x[2026];
                        n_Body_y[2027] = c_Body_y[2026];
                    end else begin
                        n_Body_x[2027] = c_Body_x[c_Size-1];
                        n_Body_y[2027] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2028) begin
                        n_Body_x[2028] = c_Body_x[2027];
                        n_Body_y[2028] = c_Body_y[2027];
                    end else begin
                        n_Body_x[2028] = c_Body_x[c_Size-1];
                        n_Body_y[2028] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2029) begin
                        n_Body_x[2029] = c_Body_x[2028];
                        n_Body_y[2029] = c_Body_y[2028];
                    end else begin
                        n_Body_x[2029] = c_Body_x[c_Size-1];
                        n_Body_y[2029] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2030) begin
                        n_Body_x[2030] = c_Body_x[2029];
                        n_Body_y[2030] = c_Body_y[2029];
                    end else begin
                        n_Body_x[2030] = c_Body_x[c_Size-1];
                        n_Body_y[2030] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2031) begin
                        n_Body_x[2031] = c_Body_x[2030];
                        n_Body_y[2031] = c_Body_y[2030];
                    end else begin
                        n_Body_x[2031] = c_Body_x[c_Size-1];
                        n_Body_y[2031] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2032) begin
                        n_Body_x[2032] = c_Body_x[2031];
                        n_Body_y[2032] = c_Body_y[2031];
                    end else begin
                        n_Body_x[2032] = c_Body_x[c_Size-1];
                        n_Body_y[2032] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2033) begin
                        n_Body_x[2033] = c_Body_x[2032];
                        n_Body_y[2033] = c_Body_y[2032];
                    end else begin
                        n_Body_x[2033] = c_Body_x[c_Size-1];
                        n_Body_y[2033] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2034) begin
                        n_Body_x[2034] = c_Body_x[2033];
                        n_Body_y[2034] = c_Body_y[2033];
                    end else begin
                        n_Body_x[2034] = c_Body_x[c_Size-1];
                        n_Body_y[2034] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2035) begin
                        n_Body_x[2035] = c_Body_x[2034];
                        n_Body_y[2035] = c_Body_y[2034];
                    end else begin
                        n_Body_x[2035] = c_Body_x[c_Size-1];
                        n_Body_y[2035] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2036) begin
                        n_Body_x[2036] = c_Body_x[2035];
                        n_Body_y[2036] = c_Body_y[2035];
                    end else begin
                        n_Body_x[2036] = c_Body_x[c_Size-1];
                        n_Body_y[2036] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2037) begin
                        n_Body_x[2037] = c_Body_x[2036];
                        n_Body_y[2037] = c_Body_y[2036];
                    end else begin
                        n_Body_x[2037] = c_Body_x[c_Size-1];
                        n_Body_y[2037] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2038) begin
                        n_Body_x[2038] = c_Body_x[2037];
                        n_Body_y[2038] = c_Body_y[2037];
                    end else begin
                        n_Body_x[2038] = c_Body_x[c_Size-1];
                        n_Body_y[2038] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2039) begin
                        n_Body_x[2039] = c_Body_x[2038];
                        n_Body_y[2039] = c_Body_y[2038];
                    end else begin
                        n_Body_x[2039] = c_Body_x[c_Size-1];
                        n_Body_y[2039] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2040) begin
                        n_Body_x[2040] = c_Body_x[2039];
                        n_Body_y[2040] = c_Body_y[2039];
                    end else begin
                        n_Body_x[2040] = c_Body_x[c_Size-1];
                        n_Body_y[2040] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2041) begin
                        n_Body_x[2041] = c_Body_x[2040];
                        n_Body_y[2041] = c_Body_y[2040];
                    end else begin
                        n_Body_x[2041] = c_Body_x[c_Size-1];
                        n_Body_y[2041] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2042) begin
                        n_Body_x[2042] = c_Body_x[2041];
                        n_Body_y[2042] = c_Body_y[2041];
                    end else begin
                        n_Body_x[2042] = c_Body_x[c_Size-1];
                        n_Body_y[2042] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2043) begin
                        n_Body_x[2043] = c_Body_x[2042];
                        n_Body_y[2043] = c_Body_y[2042];
                    end else begin
                        n_Body_x[2043] = c_Body_x[c_Size-1];
                        n_Body_y[2043] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2044) begin
                        n_Body_x[2044] = c_Body_x[2043];
                        n_Body_y[2044] = c_Body_y[2043];
                    end else begin
                        n_Body_x[2044] = c_Body_x[c_Size-1];
                        n_Body_y[2044] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2045) begin
                        n_Body_x[2045] = c_Body_x[2044];
                        n_Body_y[2045] = c_Body_y[2044];
                    end else begin
                        n_Body_x[2045] = c_Body_x[c_Size-1];
                        n_Body_y[2045] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2046) begin
                        n_Body_x[2046] = c_Body_x[2045];
                        n_Body_y[2046] = c_Body_y[2045];
                    end else begin
                        n_Body_x[2046] = c_Body_x[c_Size-1];
                        n_Body_y[2046] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2047) begin
                        n_Body_x[2047] = c_Body_x[2046];
                        n_Body_y[2047] = c_Body_y[2046];
                    end else begin
                        n_Body_x[2047] = c_Body_x[c_Size-1];
                        n_Body_y[2047] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2048) begin
                        n_Body_x[2048] = c_Body_x[2047];
                        n_Body_y[2048] = c_Body_y[2047];
                    end else begin
                        n_Body_x[2048] = c_Body_x[c_Size-1];
                        n_Body_y[2048] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2049) begin
                        n_Body_x[2049] = c_Body_x[2048];
                        n_Body_y[2049] = c_Body_y[2048];
                    end else begin
                        n_Body_x[2049] = c_Body_x[c_Size-1];
                        n_Body_y[2049] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2050) begin
                        n_Body_x[2050] = c_Body_x[2049];
                        n_Body_y[2050] = c_Body_y[2049];
                    end else begin
                        n_Body_x[2050] = c_Body_x[c_Size-1];
                        n_Body_y[2050] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2051) begin
                        n_Body_x[2051] = c_Body_x[2050];
                        n_Body_y[2051] = c_Body_y[2050];
                    end else begin
                        n_Body_x[2051] = c_Body_x[c_Size-1];
                        n_Body_y[2051] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2052) begin
                        n_Body_x[2052] = c_Body_x[2051];
                        n_Body_y[2052] = c_Body_y[2051];
                    end else begin
                        n_Body_x[2052] = c_Body_x[c_Size-1];
                        n_Body_y[2052] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2053) begin
                        n_Body_x[2053] = c_Body_x[2052];
                        n_Body_y[2053] = c_Body_y[2052];
                    end else begin
                        n_Body_x[2053] = c_Body_x[c_Size-1];
                        n_Body_y[2053] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2054) begin
                        n_Body_x[2054] = c_Body_x[2053];
                        n_Body_y[2054] = c_Body_y[2053];
                    end else begin
                        n_Body_x[2054] = c_Body_x[c_Size-1];
                        n_Body_y[2054] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2055) begin
                        n_Body_x[2055] = c_Body_x[2054];
                        n_Body_y[2055] = c_Body_y[2054];
                    end else begin
                        n_Body_x[2055] = c_Body_x[c_Size-1];
                        n_Body_y[2055] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2056) begin
                        n_Body_x[2056] = c_Body_x[2055];
                        n_Body_y[2056] = c_Body_y[2055];
                    end else begin
                        n_Body_x[2056] = c_Body_x[c_Size-1];
                        n_Body_y[2056] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2057) begin
                        n_Body_x[2057] = c_Body_x[2056];
                        n_Body_y[2057] = c_Body_y[2056];
                    end else begin
                        n_Body_x[2057] = c_Body_x[c_Size-1];
                        n_Body_y[2057] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2058) begin
                        n_Body_x[2058] = c_Body_x[2057];
                        n_Body_y[2058] = c_Body_y[2057];
                    end else begin
                        n_Body_x[2058] = c_Body_x[c_Size-1];
                        n_Body_y[2058] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2059) begin
                        n_Body_x[2059] = c_Body_x[2058];
                        n_Body_y[2059] = c_Body_y[2058];
                    end else begin
                        n_Body_x[2059] = c_Body_x[c_Size-1];
                        n_Body_y[2059] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2060) begin
                        n_Body_x[2060] = c_Body_x[2059];
                        n_Body_y[2060] = c_Body_y[2059];
                    end else begin
                        n_Body_x[2060] = c_Body_x[c_Size-1];
                        n_Body_y[2060] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2061) begin
                        n_Body_x[2061] = c_Body_x[2060];
                        n_Body_y[2061] = c_Body_y[2060];
                    end else begin
                        n_Body_x[2061] = c_Body_x[c_Size-1];
                        n_Body_y[2061] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2062) begin
                        n_Body_x[2062] = c_Body_x[2061];
                        n_Body_y[2062] = c_Body_y[2061];
                    end else begin
                        n_Body_x[2062] = c_Body_x[c_Size-1];
                        n_Body_y[2062] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2063) begin
                        n_Body_x[2063] = c_Body_x[2062];
                        n_Body_y[2063] = c_Body_y[2062];
                    end else begin
                        n_Body_x[2063] = c_Body_x[c_Size-1];
                        n_Body_y[2063] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2064) begin
                        n_Body_x[2064] = c_Body_x[2063];
                        n_Body_y[2064] = c_Body_y[2063];
                    end else begin
                        n_Body_x[2064] = c_Body_x[c_Size-1];
                        n_Body_y[2064] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2065) begin
                        n_Body_x[2065] = c_Body_x[2064];
                        n_Body_y[2065] = c_Body_y[2064];
                    end else begin
                        n_Body_x[2065] = c_Body_x[c_Size-1];
                        n_Body_y[2065] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2066) begin
                        n_Body_x[2066] = c_Body_x[2065];
                        n_Body_y[2066] = c_Body_y[2065];
                    end else begin
                        n_Body_x[2066] = c_Body_x[c_Size-1];
                        n_Body_y[2066] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2067) begin
                        n_Body_x[2067] = c_Body_x[2066];
                        n_Body_y[2067] = c_Body_y[2066];
                    end else begin
                        n_Body_x[2067] = c_Body_x[c_Size-1];
                        n_Body_y[2067] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2068) begin
                        n_Body_x[2068] = c_Body_x[2067];
                        n_Body_y[2068] = c_Body_y[2067];
                    end else begin
                        n_Body_x[2068] = c_Body_x[c_Size-1];
                        n_Body_y[2068] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2069) begin
                        n_Body_x[2069] = c_Body_x[2068];
                        n_Body_y[2069] = c_Body_y[2068];
                    end else begin
                        n_Body_x[2069] = c_Body_x[c_Size-1];
                        n_Body_y[2069] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2070) begin
                        n_Body_x[2070] = c_Body_x[2069];
                        n_Body_y[2070] = c_Body_y[2069];
                    end else begin
                        n_Body_x[2070] = c_Body_x[c_Size-1];
                        n_Body_y[2070] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2071) begin
                        n_Body_x[2071] = c_Body_x[2070];
                        n_Body_y[2071] = c_Body_y[2070];
                    end else begin
                        n_Body_x[2071] = c_Body_x[c_Size-1];
                        n_Body_y[2071] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2072) begin
                        n_Body_x[2072] = c_Body_x[2071];
                        n_Body_y[2072] = c_Body_y[2071];
                    end else begin
                        n_Body_x[2072] = c_Body_x[c_Size-1];
                        n_Body_y[2072] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2073) begin
                        n_Body_x[2073] = c_Body_x[2072];
                        n_Body_y[2073] = c_Body_y[2072];
                    end else begin
                        n_Body_x[2073] = c_Body_x[c_Size-1];
                        n_Body_y[2073] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2074) begin
                        n_Body_x[2074] = c_Body_x[2073];
                        n_Body_y[2074] = c_Body_y[2073];
                    end else begin
                        n_Body_x[2074] = c_Body_x[c_Size-1];
                        n_Body_y[2074] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2075) begin
                        n_Body_x[2075] = c_Body_x[2074];
                        n_Body_y[2075] = c_Body_y[2074];
                    end else begin
                        n_Body_x[2075] = c_Body_x[c_Size-1];
                        n_Body_y[2075] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2076) begin
                        n_Body_x[2076] = c_Body_x[2075];
                        n_Body_y[2076] = c_Body_y[2075];
                    end else begin
                        n_Body_x[2076] = c_Body_x[c_Size-1];
                        n_Body_y[2076] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2077) begin
                        n_Body_x[2077] = c_Body_x[2076];
                        n_Body_y[2077] = c_Body_y[2076];
                    end else begin
                        n_Body_x[2077] = c_Body_x[c_Size-1];
                        n_Body_y[2077] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2078) begin
                        n_Body_x[2078] = c_Body_x[2077];
                        n_Body_y[2078] = c_Body_y[2077];
                    end else begin
                        n_Body_x[2078] = c_Body_x[c_Size-1];
                        n_Body_y[2078] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2079) begin
                        n_Body_x[2079] = c_Body_x[2078];
                        n_Body_y[2079] = c_Body_y[2078];
                    end else begin
                        n_Body_x[2079] = c_Body_x[c_Size-1];
                        n_Body_y[2079] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2080) begin
                        n_Body_x[2080] = c_Body_x[2079];
                        n_Body_y[2080] = c_Body_y[2079];
                    end else begin
                        n_Body_x[2080] = c_Body_x[c_Size-1];
                        n_Body_y[2080] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2081) begin
                        n_Body_x[2081] = c_Body_x[2080];
                        n_Body_y[2081] = c_Body_y[2080];
                    end else begin
                        n_Body_x[2081] = c_Body_x[c_Size-1];
                        n_Body_y[2081] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2082) begin
                        n_Body_x[2082] = c_Body_x[2081];
                        n_Body_y[2082] = c_Body_y[2081];
                    end else begin
                        n_Body_x[2082] = c_Body_x[c_Size-1];
                        n_Body_y[2082] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2083) begin
                        n_Body_x[2083] = c_Body_x[2082];
                        n_Body_y[2083] = c_Body_y[2082];
                    end else begin
                        n_Body_x[2083] = c_Body_x[c_Size-1];
                        n_Body_y[2083] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2084) begin
                        n_Body_x[2084] = c_Body_x[2083];
                        n_Body_y[2084] = c_Body_y[2083];
                    end else begin
                        n_Body_x[2084] = c_Body_x[c_Size-1];
                        n_Body_y[2084] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2085) begin
                        n_Body_x[2085] = c_Body_x[2084];
                        n_Body_y[2085] = c_Body_y[2084];
                    end else begin
                        n_Body_x[2085] = c_Body_x[c_Size-1];
                        n_Body_y[2085] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2086) begin
                        n_Body_x[2086] = c_Body_x[2085];
                        n_Body_y[2086] = c_Body_y[2085];
                    end else begin
                        n_Body_x[2086] = c_Body_x[c_Size-1];
                        n_Body_y[2086] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2087) begin
                        n_Body_x[2087] = c_Body_x[2086];
                        n_Body_y[2087] = c_Body_y[2086];
                    end else begin
                        n_Body_x[2087] = c_Body_x[c_Size-1];
                        n_Body_y[2087] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2088) begin
                        n_Body_x[2088] = c_Body_x[2087];
                        n_Body_y[2088] = c_Body_y[2087];
                    end else begin
                        n_Body_x[2088] = c_Body_x[c_Size-1];
                        n_Body_y[2088] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2089) begin
                        n_Body_x[2089] = c_Body_x[2088];
                        n_Body_y[2089] = c_Body_y[2088];
                    end else begin
                        n_Body_x[2089] = c_Body_x[c_Size-1];
                        n_Body_y[2089] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2090) begin
                        n_Body_x[2090] = c_Body_x[2089];
                        n_Body_y[2090] = c_Body_y[2089];
                    end else begin
                        n_Body_x[2090] = c_Body_x[c_Size-1];
                        n_Body_y[2090] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2091) begin
                        n_Body_x[2091] = c_Body_x[2090];
                        n_Body_y[2091] = c_Body_y[2090];
                    end else begin
                        n_Body_x[2091] = c_Body_x[c_Size-1];
                        n_Body_y[2091] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2092) begin
                        n_Body_x[2092] = c_Body_x[2091];
                        n_Body_y[2092] = c_Body_y[2091];
                    end else begin
                        n_Body_x[2092] = c_Body_x[c_Size-1];
                        n_Body_y[2092] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2093) begin
                        n_Body_x[2093] = c_Body_x[2092];
                        n_Body_y[2093] = c_Body_y[2092];
                    end else begin
                        n_Body_x[2093] = c_Body_x[c_Size-1];
                        n_Body_y[2093] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2094) begin
                        n_Body_x[2094] = c_Body_x[2093];
                        n_Body_y[2094] = c_Body_y[2093];
                    end else begin
                        n_Body_x[2094] = c_Body_x[c_Size-1];
                        n_Body_y[2094] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2095) begin
                        n_Body_x[2095] = c_Body_x[2094];
                        n_Body_y[2095] = c_Body_y[2094];
                    end else begin
                        n_Body_x[2095] = c_Body_x[c_Size-1];
                        n_Body_y[2095] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2096) begin
                        n_Body_x[2096] = c_Body_x[2095];
                        n_Body_y[2096] = c_Body_y[2095];
                    end else begin
                        n_Body_x[2096] = c_Body_x[c_Size-1];
                        n_Body_y[2096] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2097) begin
                        n_Body_x[2097] = c_Body_x[2096];
                        n_Body_y[2097] = c_Body_y[2096];
                    end else begin
                        n_Body_x[2097] = c_Body_x[c_Size-1];
                        n_Body_y[2097] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2098) begin
                        n_Body_x[2098] = c_Body_x[2097];
                        n_Body_y[2098] = c_Body_y[2097];
                    end else begin
                        n_Body_x[2098] = c_Body_x[c_Size-1];
                        n_Body_y[2098] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2099) begin
                        n_Body_x[2099] = c_Body_x[2098];
                        n_Body_y[2099] = c_Body_y[2098];
                    end else begin
                        n_Body_x[2099] = c_Body_x[c_Size-1];
                        n_Body_y[2099] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2100) begin
                        n_Body_x[2100] = c_Body_x[2099];
                        n_Body_y[2100] = c_Body_y[2099];
                    end else begin
                        n_Body_x[2100] = c_Body_x[c_Size-1];
                        n_Body_y[2100] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2101) begin
                        n_Body_x[2101] = c_Body_x[2100];
                        n_Body_y[2101] = c_Body_y[2100];
                    end else begin
                        n_Body_x[2101] = c_Body_x[c_Size-1];
                        n_Body_y[2101] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2102) begin
                        n_Body_x[2102] = c_Body_x[2101];
                        n_Body_y[2102] = c_Body_y[2101];
                    end else begin
                        n_Body_x[2102] = c_Body_x[c_Size-1];
                        n_Body_y[2102] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2103) begin
                        n_Body_x[2103] = c_Body_x[2102];
                        n_Body_y[2103] = c_Body_y[2102];
                    end else begin
                        n_Body_x[2103] = c_Body_x[c_Size-1];
                        n_Body_y[2103] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2104) begin
                        n_Body_x[2104] = c_Body_x[2103];
                        n_Body_y[2104] = c_Body_y[2103];
                    end else begin
                        n_Body_x[2104] = c_Body_x[c_Size-1];
                        n_Body_y[2104] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2105) begin
                        n_Body_x[2105] = c_Body_x[2104];
                        n_Body_y[2105] = c_Body_y[2104];
                    end else begin
                        n_Body_x[2105] = c_Body_x[c_Size-1];
                        n_Body_y[2105] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2106) begin
                        n_Body_x[2106] = c_Body_x[2105];
                        n_Body_y[2106] = c_Body_y[2105];
                    end else begin
                        n_Body_x[2106] = c_Body_x[c_Size-1];
                        n_Body_y[2106] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2107) begin
                        n_Body_x[2107] = c_Body_x[2106];
                        n_Body_y[2107] = c_Body_y[2106];
                    end else begin
                        n_Body_x[2107] = c_Body_x[c_Size-1];
                        n_Body_y[2107] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2108) begin
                        n_Body_x[2108] = c_Body_x[2107];
                        n_Body_y[2108] = c_Body_y[2107];
                    end else begin
                        n_Body_x[2108] = c_Body_x[c_Size-1];
                        n_Body_y[2108] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2109) begin
                        n_Body_x[2109] = c_Body_x[2108];
                        n_Body_y[2109] = c_Body_y[2108];
                    end else begin
                        n_Body_x[2109] = c_Body_x[c_Size-1];
                        n_Body_y[2109] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2110) begin
                        n_Body_x[2110] = c_Body_x[2109];
                        n_Body_y[2110] = c_Body_y[2109];
                    end else begin
                        n_Body_x[2110] = c_Body_x[c_Size-1];
                        n_Body_y[2110] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2111) begin
                        n_Body_x[2111] = c_Body_x[2110];
                        n_Body_y[2111] = c_Body_y[2110];
                    end else begin
                        n_Body_x[2111] = c_Body_x[c_Size-1];
                        n_Body_y[2111] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2112) begin
                        n_Body_x[2112] = c_Body_x[2111];
                        n_Body_y[2112] = c_Body_y[2111];
                    end else begin
                        n_Body_x[2112] = c_Body_x[c_Size-1];
                        n_Body_y[2112] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2113) begin
                        n_Body_x[2113] = c_Body_x[2112];
                        n_Body_y[2113] = c_Body_y[2112];
                    end else begin
                        n_Body_x[2113] = c_Body_x[c_Size-1];
                        n_Body_y[2113] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2114) begin
                        n_Body_x[2114] = c_Body_x[2113];
                        n_Body_y[2114] = c_Body_y[2113];
                    end else begin
                        n_Body_x[2114] = c_Body_x[c_Size-1];
                        n_Body_y[2114] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2115) begin
                        n_Body_x[2115] = c_Body_x[2114];
                        n_Body_y[2115] = c_Body_y[2114];
                    end else begin
                        n_Body_x[2115] = c_Body_x[c_Size-1];
                        n_Body_y[2115] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2116) begin
                        n_Body_x[2116] = c_Body_x[2115];
                        n_Body_y[2116] = c_Body_y[2115];
                    end else begin
                        n_Body_x[2116] = c_Body_x[c_Size-1];
                        n_Body_y[2116] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2117) begin
                        n_Body_x[2117] = c_Body_x[2116];
                        n_Body_y[2117] = c_Body_y[2116];
                    end else begin
                        n_Body_x[2117] = c_Body_x[c_Size-1];
                        n_Body_y[2117] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2118) begin
                        n_Body_x[2118] = c_Body_x[2117];
                        n_Body_y[2118] = c_Body_y[2117];
                    end else begin
                        n_Body_x[2118] = c_Body_x[c_Size-1];
                        n_Body_y[2118] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2119) begin
                        n_Body_x[2119] = c_Body_x[2118];
                        n_Body_y[2119] = c_Body_y[2118];
                    end else begin
                        n_Body_x[2119] = c_Body_x[c_Size-1];
                        n_Body_y[2119] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2120) begin
                        n_Body_x[2120] = c_Body_x[2119];
                        n_Body_y[2120] = c_Body_y[2119];
                    end else begin
                        n_Body_x[2120] = c_Body_x[c_Size-1];
                        n_Body_y[2120] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2121) begin
                        n_Body_x[2121] = c_Body_x[2120];
                        n_Body_y[2121] = c_Body_y[2120];
                    end else begin
                        n_Body_x[2121] = c_Body_x[c_Size-1];
                        n_Body_y[2121] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2122) begin
                        n_Body_x[2122] = c_Body_x[2121];
                        n_Body_y[2122] = c_Body_y[2121];
                    end else begin
                        n_Body_x[2122] = c_Body_x[c_Size-1];
                        n_Body_y[2122] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2123) begin
                        n_Body_x[2123] = c_Body_x[2122];
                        n_Body_y[2123] = c_Body_y[2122];
                    end else begin
                        n_Body_x[2123] = c_Body_x[c_Size-1];
                        n_Body_y[2123] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2124) begin
                        n_Body_x[2124] = c_Body_x[2123];
                        n_Body_y[2124] = c_Body_y[2123];
                    end else begin
                        n_Body_x[2124] = c_Body_x[c_Size-1];
                        n_Body_y[2124] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2125) begin
                        n_Body_x[2125] = c_Body_x[2124];
                        n_Body_y[2125] = c_Body_y[2124];
                    end else begin
                        n_Body_x[2125] = c_Body_x[c_Size-1];
                        n_Body_y[2125] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2126) begin
                        n_Body_x[2126] = c_Body_x[2125];
                        n_Body_y[2126] = c_Body_y[2125];
                    end else begin
                        n_Body_x[2126] = c_Body_x[c_Size-1];
                        n_Body_y[2126] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2127) begin
                        n_Body_x[2127] = c_Body_x[2126];
                        n_Body_y[2127] = c_Body_y[2126];
                    end else begin
                        n_Body_x[2127] = c_Body_x[c_Size-1];
                        n_Body_y[2127] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2128) begin
                        n_Body_x[2128] = c_Body_x[2127];
                        n_Body_y[2128] = c_Body_y[2127];
                    end else begin
                        n_Body_x[2128] = c_Body_x[c_Size-1];
                        n_Body_y[2128] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2129) begin
                        n_Body_x[2129] = c_Body_x[2128];
                        n_Body_y[2129] = c_Body_y[2128];
                    end else begin
                        n_Body_x[2129] = c_Body_x[c_Size-1];
                        n_Body_y[2129] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2130) begin
                        n_Body_x[2130] = c_Body_x[2129];
                        n_Body_y[2130] = c_Body_y[2129];
                    end else begin
                        n_Body_x[2130] = c_Body_x[c_Size-1];
                        n_Body_y[2130] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2131) begin
                        n_Body_x[2131] = c_Body_x[2130];
                        n_Body_y[2131] = c_Body_y[2130];
                    end else begin
                        n_Body_x[2131] = c_Body_x[c_Size-1];
                        n_Body_y[2131] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2132) begin
                        n_Body_x[2132] = c_Body_x[2131];
                        n_Body_y[2132] = c_Body_y[2131];
                    end else begin
                        n_Body_x[2132] = c_Body_x[c_Size-1];
                        n_Body_y[2132] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2133) begin
                        n_Body_x[2133] = c_Body_x[2132];
                        n_Body_y[2133] = c_Body_y[2132];
                    end else begin
                        n_Body_x[2133] = c_Body_x[c_Size-1];
                        n_Body_y[2133] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2134) begin
                        n_Body_x[2134] = c_Body_x[2133];
                        n_Body_y[2134] = c_Body_y[2133];
                    end else begin
                        n_Body_x[2134] = c_Body_x[c_Size-1];
                        n_Body_y[2134] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2135) begin
                        n_Body_x[2135] = c_Body_x[2134];
                        n_Body_y[2135] = c_Body_y[2134];
                    end else begin
                        n_Body_x[2135] = c_Body_x[c_Size-1];
                        n_Body_y[2135] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2136) begin
                        n_Body_x[2136] = c_Body_x[2135];
                        n_Body_y[2136] = c_Body_y[2135];
                    end else begin
                        n_Body_x[2136] = c_Body_x[c_Size-1];
                        n_Body_y[2136] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2137) begin
                        n_Body_x[2137] = c_Body_x[2136];
                        n_Body_y[2137] = c_Body_y[2136];
                    end else begin
                        n_Body_x[2137] = c_Body_x[c_Size-1];
                        n_Body_y[2137] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2138) begin
                        n_Body_x[2138] = c_Body_x[2137];
                        n_Body_y[2138] = c_Body_y[2137];
                    end else begin
                        n_Body_x[2138] = c_Body_x[c_Size-1];
                        n_Body_y[2138] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2139) begin
                        n_Body_x[2139] = c_Body_x[2138];
                        n_Body_y[2139] = c_Body_y[2138];
                    end else begin
                        n_Body_x[2139] = c_Body_x[c_Size-1];
                        n_Body_y[2139] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2140) begin
                        n_Body_x[2140] = c_Body_x[2139];
                        n_Body_y[2140] = c_Body_y[2139];
                    end else begin
                        n_Body_x[2140] = c_Body_x[c_Size-1];
                        n_Body_y[2140] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2141) begin
                        n_Body_x[2141] = c_Body_x[2140];
                        n_Body_y[2141] = c_Body_y[2140];
                    end else begin
                        n_Body_x[2141] = c_Body_x[c_Size-1];
                        n_Body_y[2141] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2142) begin
                        n_Body_x[2142] = c_Body_x[2141];
                        n_Body_y[2142] = c_Body_y[2141];
                    end else begin
                        n_Body_x[2142] = c_Body_x[c_Size-1];
                        n_Body_y[2142] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2143) begin
                        n_Body_x[2143] = c_Body_x[2142];
                        n_Body_y[2143] = c_Body_y[2142];
                    end else begin
                        n_Body_x[2143] = c_Body_x[c_Size-1];
                        n_Body_y[2143] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2144) begin
                        n_Body_x[2144] = c_Body_x[2143];
                        n_Body_y[2144] = c_Body_y[2143];
                    end else begin
                        n_Body_x[2144] = c_Body_x[c_Size-1];
                        n_Body_y[2144] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2145) begin
                        n_Body_x[2145] = c_Body_x[2144];
                        n_Body_y[2145] = c_Body_y[2144];
                    end else begin
                        n_Body_x[2145] = c_Body_x[c_Size-1];
                        n_Body_y[2145] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2146) begin
                        n_Body_x[2146] = c_Body_x[2145];
                        n_Body_y[2146] = c_Body_y[2145];
                    end else begin
                        n_Body_x[2146] = c_Body_x[c_Size-1];
                        n_Body_y[2146] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2147) begin
                        n_Body_x[2147] = c_Body_x[2146];
                        n_Body_y[2147] = c_Body_y[2146];
                    end else begin
                        n_Body_x[2147] = c_Body_x[c_Size-1];
                        n_Body_y[2147] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2148) begin
                        n_Body_x[2148] = c_Body_x[2147];
                        n_Body_y[2148] = c_Body_y[2147];
                    end else begin
                        n_Body_x[2148] = c_Body_x[c_Size-1];
                        n_Body_y[2148] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2149) begin
                        n_Body_x[2149] = c_Body_x[2148];
                        n_Body_y[2149] = c_Body_y[2148];
                    end else begin
                        n_Body_x[2149] = c_Body_x[c_Size-1];
                        n_Body_y[2149] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2150) begin
                        n_Body_x[2150] = c_Body_x[2149];
                        n_Body_y[2150] = c_Body_y[2149];
                    end else begin
                        n_Body_x[2150] = c_Body_x[c_Size-1];
                        n_Body_y[2150] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2151) begin
                        n_Body_x[2151] = c_Body_x[2150];
                        n_Body_y[2151] = c_Body_y[2150];
                    end else begin
                        n_Body_x[2151] = c_Body_x[c_Size-1];
                        n_Body_y[2151] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2152) begin
                        n_Body_x[2152] = c_Body_x[2151];
                        n_Body_y[2152] = c_Body_y[2151];
                    end else begin
                        n_Body_x[2152] = c_Body_x[c_Size-1];
                        n_Body_y[2152] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2153) begin
                        n_Body_x[2153] = c_Body_x[2152];
                        n_Body_y[2153] = c_Body_y[2152];
                    end else begin
                        n_Body_x[2153] = c_Body_x[c_Size-1];
                        n_Body_y[2153] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2154) begin
                        n_Body_x[2154] = c_Body_x[2153];
                        n_Body_y[2154] = c_Body_y[2153];
                    end else begin
                        n_Body_x[2154] = c_Body_x[c_Size-1];
                        n_Body_y[2154] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2155) begin
                        n_Body_x[2155] = c_Body_x[2154];
                        n_Body_y[2155] = c_Body_y[2154];
                    end else begin
                        n_Body_x[2155] = c_Body_x[c_Size-1];
                        n_Body_y[2155] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2156) begin
                        n_Body_x[2156] = c_Body_x[2155];
                        n_Body_y[2156] = c_Body_y[2155];
                    end else begin
                        n_Body_x[2156] = c_Body_x[c_Size-1];
                        n_Body_y[2156] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2157) begin
                        n_Body_x[2157] = c_Body_x[2156];
                        n_Body_y[2157] = c_Body_y[2156];
                    end else begin
                        n_Body_x[2157] = c_Body_x[c_Size-1];
                        n_Body_y[2157] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2158) begin
                        n_Body_x[2158] = c_Body_x[2157];
                        n_Body_y[2158] = c_Body_y[2157];
                    end else begin
                        n_Body_x[2158] = c_Body_x[c_Size-1];
                        n_Body_y[2158] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2159) begin
                        n_Body_x[2159] = c_Body_x[2158];
                        n_Body_y[2159] = c_Body_y[2158];
                    end else begin
                        n_Body_x[2159] = c_Body_x[c_Size-1];
                        n_Body_y[2159] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2160) begin
                        n_Body_x[2160] = c_Body_x[2159];
                        n_Body_y[2160] = c_Body_y[2159];
                    end else begin
                        n_Body_x[2160] = c_Body_x[c_Size-1];
                        n_Body_y[2160] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2161) begin
                        n_Body_x[2161] = c_Body_x[2160];
                        n_Body_y[2161] = c_Body_y[2160];
                    end else begin
                        n_Body_x[2161] = c_Body_x[c_Size-1];
                        n_Body_y[2161] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2162) begin
                        n_Body_x[2162] = c_Body_x[2161];
                        n_Body_y[2162] = c_Body_y[2161];
                    end else begin
                        n_Body_x[2162] = c_Body_x[c_Size-1];
                        n_Body_y[2162] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2163) begin
                        n_Body_x[2163] = c_Body_x[2162];
                        n_Body_y[2163] = c_Body_y[2162];
                    end else begin
                        n_Body_x[2163] = c_Body_x[c_Size-1];
                        n_Body_y[2163] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2164) begin
                        n_Body_x[2164] = c_Body_x[2163];
                        n_Body_y[2164] = c_Body_y[2163];
                    end else begin
                        n_Body_x[2164] = c_Body_x[c_Size-1];
                        n_Body_y[2164] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2165) begin
                        n_Body_x[2165] = c_Body_x[2164];
                        n_Body_y[2165] = c_Body_y[2164];
                    end else begin
                        n_Body_x[2165] = c_Body_x[c_Size-1];
                        n_Body_y[2165] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2166) begin
                        n_Body_x[2166] = c_Body_x[2165];
                        n_Body_y[2166] = c_Body_y[2165];
                    end else begin
                        n_Body_x[2166] = c_Body_x[c_Size-1];
                        n_Body_y[2166] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2167) begin
                        n_Body_x[2167] = c_Body_x[2166];
                        n_Body_y[2167] = c_Body_y[2166];
                    end else begin
                        n_Body_x[2167] = c_Body_x[c_Size-1];
                        n_Body_y[2167] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2168) begin
                        n_Body_x[2168] = c_Body_x[2167];
                        n_Body_y[2168] = c_Body_y[2167];
                    end else begin
                        n_Body_x[2168] = c_Body_x[c_Size-1];
                        n_Body_y[2168] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2169) begin
                        n_Body_x[2169] = c_Body_x[2168];
                        n_Body_y[2169] = c_Body_y[2168];
                    end else begin
                        n_Body_x[2169] = c_Body_x[c_Size-1];
                        n_Body_y[2169] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2170) begin
                        n_Body_x[2170] = c_Body_x[2169];
                        n_Body_y[2170] = c_Body_y[2169];
                    end else begin
                        n_Body_x[2170] = c_Body_x[c_Size-1];
                        n_Body_y[2170] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2171) begin
                        n_Body_x[2171] = c_Body_x[2170];
                        n_Body_y[2171] = c_Body_y[2170];
                    end else begin
                        n_Body_x[2171] = c_Body_x[c_Size-1];
                        n_Body_y[2171] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2172) begin
                        n_Body_x[2172] = c_Body_x[2171];
                        n_Body_y[2172] = c_Body_y[2171];
                    end else begin
                        n_Body_x[2172] = c_Body_x[c_Size-1];
                        n_Body_y[2172] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2173) begin
                        n_Body_x[2173] = c_Body_x[2172];
                        n_Body_y[2173] = c_Body_y[2172];
                    end else begin
                        n_Body_x[2173] = c_Body_x[c_Size-1];
                        n_Body_y[2173] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2174) begin
                        n_Body_x[2174] = c_Body_x[2173];
                        n_Body_y[2174] = c_Body_y[2173];
                    end else begin
                        n_Body_x[2174] = c_Body_x[c_Size-1];
                        n_Body_y[2174] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2175) begin
                        n_Body_x[2175] = c_Body_x[2174];
                        n_Body_y[2175] = c_Body_y[2174];
                    end else begin
                        n_Body_x[2175] = c_Body_x[c_Size-1];
                        n_Body_y[2175] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2176) begin
                        n_Body_x[2176] = c_Body_x[2175];
                        n_Body_y[2176] = c_Body_y[2175];
                    end else begin
                        n_Body_x[2176] = c_Body_x[c_Size-1];
                        n_Body_y[2176] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2177) begin
                        n_Body_x[2177] = c_Body_x[2176];
                        n_Body_y[2177] = c_Body_y[2176];
                    end else begin
                        n_Body_x[2177] = c_Body_x[c_Size-1];
                        n_Body_y[2177] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2178) begin
                        n_Body_x[2178] = c_Body_x[2177];
                        n_Body_y[2178] = c_Body_y[2177];
                    end else begin
                        n_Body_x[2178] = c_Body_x[c_Size-1];
                        n_Body_y[2178] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2179) begin
                        n_Body_x[2179] = c_Body_x[2178];
                        n_Body_y[2179] = c_Body_y[2178];
                    end else begin
                        n_Body_x[2179] = c_Body_x[c_Size-1];
                        n_Body_y[2179] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2180) begin
                        n_Body_x[2180] = c_Body_x[2179];
                        n_Body_y[2180] = c_Body_y[2179];
                    end else begin
                        n_Body_x[2180] = c_Body_x[c_Size-1];
                        n_Body_y[2180] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2181) begin
                        n_Body_x[2181] = c_Body_x[2180];
                        n_Body_y[2181] = c_Body_y[2180];
                    end else begin
                        n_Body_x[2181] = c_Body_x[c_Size-1];
                        n_Body_y[2181] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2182) begin
                        n_Body_x[2182] = c_Body_x[2181];
                        n_Body_y[2182] = c_Body_y[2181];
                    end else begin
                        n_Body_x[2182] = c_Body_x[c_Size-1];
                        n_Body_y[2182] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2183) begin
                        n_Body_x[2183] = c_Body_x[2182];
                        n_Body_y[2183] = c_Body_y[2182];
                    end else begin
                        n_Body_x[2183] = c_Body_x[c_Size-1];
                        n_Body_y[2183] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2184) begin
                        n_Body_x[2184] = c_Body_x[2183];
                        n_Body_y[2184] = c_Body_y[2183];
                    end else begin
                        n_Body_x[2184] = c_Body_x[c_Size-1];
                        n_Body_y[2184] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2185) begin
                        n_Body_x[2185] = c_Body_x[2184];
                        n_Body_y[2185] = c_Body_y[2184];
                    end else begin
                        n_Body_x[2185] = c_Body_x[c_Size-1];
                        n_Body_y[2185] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2186) begin
                        n_Body_x[2186] = c_Body_x[2185];
                        n_Body_y[2186] = c_Body_y[2185];
                    end else begin
                        n_Body_x[2186] = c_Body_x[c_Size-1];
                        n_Body_y[2186] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2187) begin
                        n_Body_x[2187] = c_Body_x[2186];
                        n_Body_y[2187] = c_Body_y[2186];
                    end else begin
                        n_Body_x[2187] = c_Body_x[c_Size-1];
                        n_Body_y[2187] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2188) begin
                        n_Body_x[2188] = c_Body_x[2187];
                        n_Body_y[2188] = c_Body_y[2187];
                    end else begin
                        n_Body_x[2188] = c_Body_x[c_Size-1];
                        n_Body_y[2188] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2189) begin
                        n_Body_x[2189] = c_Body_x[2188];
                        n_Body_y[2189] = c_Body_y[2188];
                    end else begin
                        n_Body_x[2189] = c_Body_x[c_Size-1];
                        n_Body_y[2189] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2190) begin
                        n_Body_x[2190] = c_Body_x[2189];
                        n_Body_y[2190] = c_Body_y[2189];
                    end else begin
                        n_Body_x[2190] = c_Body_x[c_Size-1];
                        n_Body_y[2190] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2191) begin
                        n_Body_x[2191] = c_Body_x[2190];
                        n_Body_y[2191] = c_Body_y[2190];
                    end else begin
                        n_Body_x[2191] = c_Body_x[c_Size-1];
                        n_Body_y[2191] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2192) begin
                        n_Body_x[2192] = c_Body_x[2191];
                        n_Body_y[2192] = c_Body_y[2191];
                    end else begin
                        n_Body_x[2192] = c_Body_x[c_Size-1];
                        n_Body_y[2192] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2193) begin
                        n_Body_x[2193] = c_Body_x[2192];
                        n_Body_y[2193] = c_Body_y[2192];
                    end else begin
                        n_Body_x[2193] = c_Body_x[c_Size-1];
                        n_Body_y[2193] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2194) begin
                        n_Body_x[2194] = c_Body_x[2193];
                        n_Body_y[2194] = c_Body_y[2193];
                    end else begin
                        n_Body_x[2194] = c_Body_x[c_Size-1];
                        n_Body_y[2194] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2195) begin
                        n_Body_x[2195] = c_Body_x[2194];
                        n_Body_y[2195] = c_Body_y[2194];
                    end else begin
                        n_Body_x[2195] = c_Body_x[c_Size-1];
                        n_Body_y[2195] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2196) begin
                        n_Body_x[2196] = c_Body_x[2195];
                        n_Body_y[2196] = c_Body_y[2195];
                    end else begin
                        n_Body_x[2196] = c_Body_x[c_Size-1];
                        n_Body_y[2196] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2197) begin
                        n_Body_x[2197] = c_Body_x[2196];
                        n_Body_y[2197] = c_Body_y[2196];
                    end else begin
                        n_Body_x[2197] = c_Body_x[c_Size-1];
                        n_Body_y[2197] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2198) begin
                        n_Body_x[2198] = c_Body_x[2197];
                        n_Body_y[2198] = c_Body_y[2197];
                    end else begin
                        n_Body_x[2198] = c_Body_x[c_Size-1];
                        n_Body_y[2198] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2199) begin
                        n_Body_x[2199] = c_Body_x[2198];
                        n_Body_y[2199] = c_Body_y[2198];
                    end else begin
                        n_Body_x[2199] = c_Body_x[c_Size-1];
                        n_Body_y[2199] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2200) begin
                        n_Body_x[2200] = c_Body_x[2199];
                        n_Body_y[2200] = c_Body_y[2199];
                    end else begin
                        n_Body_x[2200] = c_Body_x[c_Size-1];
                        n_Body_y[2200] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2201) begin
                        n_Body_x[2201] = c_Body_x[2200];
                        n_Body_y[2201] = c_Body_y[2200];
                    end else begin
                        n_Body_x[2201] = c_Body_x[c_Size-1];
                        n_Body_y[2201] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2202) begin
                        n_Body_x[2202] = c_Body_x[2201];
                        n_Body_y[2202] = c_Body_y[2201];
                    end else begin
                        n_Body_x[2202] = c_Body_x[c_Size-1];
                        n_Body_y[2202] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2203) begin
                        n_Body_x[2203] = c_Body_x[2202];
                        n_Body_y[2203] = c_Body_y[2202];
                    end else begin
                        n_Body_x[2203] = c_Body_x[c_Size-1];
                        n_Body_y[2203] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2204) begin
                        n_Body_x[2204] = c_Body_x[2203];
                        n_Body_y[2204] = c_Body_y[2203];
                    end else begin
                        n_Body_x[2204] = c_Body_x[c_Size-1];
                        n_Body_y[2204] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2205) begin
                        n_Body_x[2205] = c_Body_x[2204];
                        n_Body_y[2205] = c_Body_y[2204];
                    end else begin
                        n_Body_x[2205] = c_Body_x[c_Size-1];
                        n_Body_y[2205] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2206) begin
                        n_Body_x[2206] = c_Body_x[2205];
                        n_Body_y[2206] = c_Body_y[2205];
                    end else begin
                        n_Body_x[2206] = c_Body_x[c_Size-1];
                        n_Body_y[2206] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2207) begin
                        n_Body_x[2207] = c_Body_x[2206];
                        n_Body_y[2207] = c_Body_y[2206];
                    end else begin
                        n_Body_x[2207] = c_Body_x[c_Size-1];
                        n_Body_y[2207] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2208) begin
                        n_Body_x[2208] = c_Body_x[2207];
                        n_Body_y[2208] = c_Body_y[2207];
                    end else begin
                        n_Body_x[2208] = c_Body_x[c_Size-1];
                        n_Body_y[2208] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2209) begin
                        n_Body_x[2209] = c_Body_x[2208];
                        n_Body_y[2209] = c_Body_y[2208];
                    end else begin
                        n_Body_x[2209] = c_Body_x[c_Size-1];
                        n_Body_y[2209] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2210) begin
                        n_Body_x[2210] = c_Body_x[2209];
                        n_Body_y[2210] = c_Body_y[2209];
                    end else begin
                        n_Body_x[2210] = c_Body_x[c_Size-1];
                        n_Body_y[2210] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2211) begin
                        n_Body_x[2211] = c_Body_x[2210];
                        n_Body_y[2211] = c_Body_y[2210];
                    end else begin
                        n_Body_x[2211] = c_Body_x[c_Size-1];
                        n_Body_y[2211] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2212) begin
                        n_Body_x[2212] = c_Body_x[2211];
                        n_Body_y[2212] = c_Body_y[2211];
                    end else begin
                        n_Body_x[2212] = c_Body_x[c_Size-1];
                        n_Body_y[2212] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2213) begin
                        n_Body_x[2213] = c_Body_x[2212];
                        n_Body_y[2213] = c_Body_y[2212];
                    end else begin
                        n_Body_x[2213] = c_Body_x[c_Size-1];
                        n_Body_y[2213] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2214) begin
                        n_Body_x[2214] = c_Body_x[2213];
                        n_Body_y[2214] = c_Body_y[2213];
                    end else begin
                        n_Body_x[2214] = c_Body_x[c_Size-1];
                        n_Body_y[2214] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2215) begin
                        n_Body_x[2215] = c_Body_x[2214];
                        n_Body_y[2215] = c_Body_y[2214];
                    end else begin
                        n_Body_x[2215] = c_Body_x[c_Size-1];
                        n_Body_y[2215] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2216) begin
                        n_Body_x[2216] = c_Body_x[2215];
                        n_Body_y[2216] = c_Body_y[2215];
                    end else begin
                        n_Body_x[2216] = c_Body_x[c_Size-1];
                        n_Body_y[2216] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2217) begin
                        n_Body_x[2217] = c_Body_x[2216];
                        n_Body_y[2217] = c_Body_y[2216];
                    end else begin
                        n_Body_x[2217] = c_Body_x[c_Size-1];
                        n_Body_y[2217] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2218) begin
                        n_Body_x[2218] = c_Body_x[2217];
                        n_Body_y[2218] = c_Body_y[2217];
                    end else begin
                        n_Body_x[2218] = c_Body_x[c_Size-1];
                        n_Body_y[2218] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2219) begin
                        n_Body_x[2219] = c_Body_x[2218];
                        n_Body_y[2219] = c_Body_y[2218];
                    end else begin
                        n_Body_x[2219] = c_Body_x[c_Size-1];
                        n_Body_y[2219] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2220) begin
                        n_Body_x[2220] = c_Body_x[2219];
                        n_Body_y[2220] = c_Body_y[2219];
                    end else begin
                        n_Body_x[2220] = c_Body_x[c_Size-1];
                        n_Body_y[2220] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2221) begin
                        n_Body_x[2221] = c_Body_x[2220];
                        n_Body_y[2221] = c_Body_y[2220];
                    end else begin
                        n_Body_x[2221] = c_Body_x[c_Size-1];
                        n_Body_y[2221] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2222) begin
                        n_Body_x[2222] = c_Body_x[2221];
                        n_Body_y[2222] = c_Body_y[2221];
                    end else begin
                        n_Body_x[2222] = c_Body_x[c_Size-1];
                        n_Body_y[2222] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2223) begin
                        n_Body_x[2223] = c_Body_x[2222];
                        n_Body_y[2223] = c_Body_y[2222];
                    end else begin
                        n_Body_x[2223] = c_Body_x[c_Size-1];
                        n_Body_y[2223] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2224) begin
                        n_Body_x[2224] = c_Body_x[2223];
                        n_Body_y[2224] = c_Body_y[2223];
                    end else begin
                        n_Body_x[2224] = c_Body_x[c_Size-1];
                        n_Body_y[2224] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2225) begin
                        n_Body_x[2225] = c_Body_x[2224];
                        n_Body_y[2225] = c_Body_y[2224];
                    end else begin
                        n_Body_x[2225] = c_Body_x[c_Size-1];
                        n_Body_y[2225] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2226) begin
                        n_Body_x[2226] = c_Body_x[2225];
                        n_Body_y[2226] = c_Body_y[2225];
                    end else begin
                        n_Body_x[2226] = c_Body_x[c_Size-1];
                        n_Body_y[2226] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2227) begin
                        n_Body_x[2227] = c_Body_x[2226];
                        n_Body_y[2227] = c_Body_y[2226];
                    end else begin
                        n_Body_x[2227] = c_Body_x[c_Size-1];
                        n_Body_y[2227] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2228) begin
                        n_Body_x[2228] = c_Body_x[2227];
                        n_Body_y[2228] = c_Body_y[2227];
                    end else begin
                        n_Body_x[2228] = c_Body_x[c_Size-1];
                        n_Body_y[2228] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2229) begin
                        n_Body_x[2229] = c_Body_x[2228];
                        n_Body_y[2229] = c_Body_y[2228];
                    end else begin
                        n_Body_x[2229] = c_Body_x[c_Size-1];
                        n_Body_y[2229] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2230) begin
                        n_Body_x[2230] = c_Body_x[2229];
                        n_Body_y[2230] = c_Body_y[2229];
                    end else begin
                        n_Body_x[2230] = c_Body_x[c_Size-1];
                        n_Body_y[2230] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2231) begin
                        n_Body_x[2231] = c_Body_x[2230];
                        n_Body_y[2231] = c_Body_y[2230];
                    end else begin
                        n_Body_x[2231] = c_Body_x[c_Size-1];
                        n_Body_y[2231] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2232) begin
                        n_Body_x[2232] = c_Body_x[2231];
                        n_Body_y[2232] = c_Body_y[2231];
                    end else begin
                        n_Body_x[2232] = c_Body_x[c_Size-1];
                        n_Body_y[2232] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2233) begin
                        n_Body_x[2233] = c_Body_x[2232];
                        n_Body_y[2233] = c_Body_y[2232];
                    end else begin
                        n_Body_x[2233] = c_Body_x[c_Size-1];
                        n_Body_y[2233] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2234) begin
                        n_Body_x[2234] = c_Body_x[2233];
                        n_Body_y[2234] = c_Body_y[2233];
                    end else begin
                        n_Body_x[2234] = c_Body_x[c_Size-1];
                        n_Body_y[2234] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2235) begin
                        n_Body_x[2235] = c_Body_x[2234];
                        n_Body_y[2235] = c_Body_y[2234];
                    end else begin
                        n_Body_x[2235] = c_Body_x[c_Size-1];
                        n_Body_y[2235] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2236) begin
                        n_Body_x[2236] = c_Body_x[2235];
                        n_Body_y[2236] = c_Body_y[2235];
                    end else begin
                        n_Body_x[2236] = c_Body_x[c_Size-1];
                        n_Body_y[2236] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2237) begin
                        n_Body_x[2237] = c_Body_x[2236];
                        n_Body_y[2237] = c_Body_y[2236];
                    end else begin
                        n_Body_x[2237] = c_Body_x[c_Size-1];
                        n_Body_y[2237] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2238) begin
                        n_Body_x[2238] = c_Body_x[2237];
                        n_Body_y[2238] = c_Body_y[2237];
                    end else begin
                        n_Body_x[2238] = c_Body_x[c_Size-1];
                        n_Body_y[2238] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2239) begin
                        n_Body_x[2239] = c_Body_x[2238];
                        n_Body_y[2239] = c_Body_y[2238];
                    end else begin
                        n_Body_x[2239] = c_Body_x[c_Size-1];
                        n_Body_y[2239] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2240) begin
                        n_Body_x[2240] = c_Body_x[2239];
                        n_Body_y[2240] = c_Body_y[2239];
                    end else begin
                        n_Body_x[2240] = c_Body_x[c_Size-1];
                        n_Body_y[2240] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2241) begin
                        n_Body_x[2241] = c_Body_x[2240];
                        n_Body_y[2241] = c_Body_y[2240];
                    end else begin
                        n_Body_x[2241] = c_Body_x[c_Size-1];
                        n_Body_y[2241] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2242) begin
                        n_Body_x[2242] = c_Body_x[2241];
                        n_Body_y[2242] = c_Body_y[2241];
                    end else begin
                        n_Body_x[2242] = c_Body_x[c_Size-1];
                        n_Body_y[2242] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2243) begin
                        n_Body_x[2243] = c_Body_x[2242];
                        n_Body_y[2243] = c_Body_y[2242];
                    end else begin
                        n_Body_x[2243] = c_Body_x[c_Size-1];
                        n_Body_y[2243] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2244) begin
                        n_Body_x[2244] = c_Body_x[2243];
                        n_Body_y[2244] = c_Body_y[2243];
                    end else begin
                        n_Body_x[2244] = c_Body_x[c_Size-1];
                        n_Body_y[2244] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2245) begin
                        n_Body_x[2245] = c_Body_x[2244];
                        n_Body_y[2245] = c_Body_y[2244];
                    end else begin
                        n_Body_x[2245] = c_Body_x[c_Size-1];
                        n_Body_y[2245] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2246) begin
                        n_Body_x[2246] = c_Body_x[2245];
                        n_Body_y[2246] = c_Body_y[2245];
                    end else begin
                        n_Body_x[2246] = c_Body_x[c_Size-1];
                        n_Body_y[2246] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2247) begin
                        n_Body_x[2247] = c_Body_x[2246];
                        n_Body_y[2247] = c_Body_y[2246];
                    end else begin
                        n_Body_x[2247] = c_Body_x[c_Size-1];
                        n_Body_y[2247] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2248) begin
                        n_Body_x[2248] = c_Body_x[2247];
                        n_Body_y[2248] = c_Body_y[2247];
                    end else begin
                        n_Body_x[2248] = c_Body_x[c_Size-1];
                        n_Body_y[2248] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2249) begin
                        n_Body_x[2249] = c_Body_x[2248];
                        n_Body_y[2249] = c_Body_y[2248];
                    end else begin
                        n_Body_x[2249] = c_Body_x[c_Size-1];
                        n_Body_y[2249] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2250) begin
                        n_Body_x[2250] = c_Body_x[2249];
                        n_Body_y[2250] = c_Body_y[2249];
                    end else begin
                        n_Body_x[2250] = c_Body_x[c_Size-1];
                        n_Body_y[2250] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2251) begin
                        n_Body_x[2251] = c_Body_x[2250];
                        n_Body_y[2251] = c_Body_y[2250];
                    end else begin
                        n_Body_x[2251] = c_Body_x[c_Size-1];
                        n_Body_y[2251] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2252) begin
                        n_Body_x[2252] = c_Body_x[2251];
                        n_Body_y[2252] = c_Body_y[2251];
                    end else begin
                        n_Body_x[2252] = c_Body_x[c_Size-1];
                        n_Body_y[2252] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2253) begin
                        n_Body_x[2253] = c_Body_x[2252];
                        n_Body_y[2253] = c_Body_y[2252];
                    end else begin
                        n_Body_x[2253] = c_Body_x[c_Size-1];
                        n_Body_y[2253] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2254) begin
                        n_Body_x[2254] = c_Body_x[2253];
                        n_Body_y[2254] = c_Body_y[2253];
                    end else begin
                        n_Body_x[2254] = c_Body_x[c_Size-1];
                        n_Body_y[2254] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2255) begin
                        n_Body_x[2255] = c_Body_x[2254];
                        n_Body_y[2255] = c_Body_y[2254];
                    end else begin
                        n_Body_x[2255] = c_Body_x[c_Size-1];
                        n_Body_y[2255] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2256) begin
                        n_Body_x[2256] = c_Body_x[2255];
                        n_Body_y[2256] = c_Body_y[2255];
                    end else begin
                        n_Body_x[2256] = c_Body_x[c_Size-1];
                        n_Body_y[2256] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2257) begin
                        n_Body_x[2257] = c_Body_x[2256];
                        n_Body_y[2257] = c_Body_y[2256];
                    end else begin
                        n_Body_x[2257] = c_Body_x[c_Size-1];
                        n_Body_y[2257] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2258) begin
                        n_Body_x[2258] = c_Body_x[2257];
                        n_Body_y[2258] = c_Body_y[2257];
                    end else begin
                        n_Body_x[2258] = c_Body_x[c_Size-1];
                        n_Body_y[2258] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2259) begin
                        n_Body_x[2259] = c_Body_x[2258];
                        n_Body_y[2259] = c_Body_y[2258];
                    end else begin
                        n_Body_x[2259] = c_Body_x[c_Size-1];
                        n_Body_y[2259] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2260) begin
                        n_Body_x[2260] = c_Body_x[2259];
                        n_Body_y[2260] = c_Body_y[2259];
                    end else begin
                        n_Body_x[2260] = c_Body_x[c_Size-1];
                        n_Body_y[2260] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2261) begin
                        n_Body_x[2261] = c_Body_x[2260];
                        n_Body_y[2261] = c_Body_y[2260];
                    end else begin
                        n_Body_x[2261] = c_Body_x[c_Size-1];
                        n_Body_y[2261] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2262) begin
                        n_Body_x[2262] = c_Body_x[2261];
                        n_Body_y[2262] = c_Body_y[2261];
                    end else begin
                        n_Body_x[2262] = c_Body_x[c_Size-1];
                        n_Body_y[2262] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2263) begin
                        n_Body_x[2263] = c_Body_x[2262];
                        n_Body_y[2263] = c_Body_y[2262];
                    end else begin
                        n_Body_x[2263] = c_Body_x[c_Size-1];
                        n_Body_y[2263] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2264) begin
                        n_Body_x[2264] = c_Body_x[2263];
                        n_Body_y[2264] = c_Body_y[2263];
                    end else begin
                        n_Body_x[2264] = c_Body_x[c_Size-1];
                        n_Body_y[2264] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2265) begin
                        n_Body_x[2265] = c_Body_x[2264];
                        n_Body_y[2265] = c_Body_y[2264];
                    end else begin
                        n_Body_x[2265] = c_Body_x[c_Size-1];
                        n_Body_y[2265] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2266) begin
                        n_Body_x[2266] = c_Body_x[2265];
                        n_Body_y[2266] = c_Body_y[2265];
                    end else begin
                        n_Body_x[2266] = c_Body_x[c_Size-1];
                        n_Body_y[2266] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2267) begin
                        n_Body_x[2267] = c_Body_x[2266];
                        n_Body_y[2267] = c_Body_y[2266];
                    end else begin
                        n_Body_x[2267] = c_Body_x[c_Size-1];
                        n_Body_y[2267] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2268) begin
                        n_Body_x[2268] = c_Body_x[2267];
                        n_Body_y[2268] = c_Body_y[2267];
                    end else begin
                        n_Body_x[2268] = c_Body_x[c_Size-1];
                        n_Body_y[2268] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2269) begin
                        n_Body_x[2269] = c_Body_x[2268];
                        n_Body_y[2269] = c_Body_y[2268];
                    end else begin
                        n_Body_x[2269] = c_Body_x[c_Size-1];
                        n_Body_y[2269] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2270) begin
                        n_Body_x[2270] = c_Body_x[2269];
                        n_Body_y[2270] = c_Body_y[2269];
                    end else begin
                        n_Body_x[2270] = c_Body_x[c_Size-1];
                        n_Body_y[2270] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2271) begin
                        n_Body_x[2271] = c_Body_x[2270];
                        n_Body_y[2271] = c_Body_y[2270];
                    end else begin
                        n_Body_x[2271] = c_Body_x[c_Size-1];
                        n_Body_y[2271] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2272) begin
                        n_Body_x[2272] = c_Body_x[2271];
                        n_Body_y[2272] = c_Body_y[2271];
                    end else begin
                        n_Body_x[2272] = c_Body_x[c_Size-1];
                        n_Body_y[2272] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2273) begin
                        n_Body_x[2273] = c_Body_x[2272];
                        n_Body_y[2273] = c_Body_y[2272];
                    end else begin
                        n_Body_x[2273] = c_Body_x[c_Size-1];
                        n_Body_y[2273] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2274) begin
                        n_Body_x[2274] = c_Body_x[2273];
                        n_Body_y[2274] = c_Body_y[2273];
                    end else begin
                        n_Body_x[2274] = c_Body_x[c_Size-1];
                        n_Body_y[2274] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2275) begin
                        n_Body_x[2275] = c_Body_x[2274];
                        n_Body_y[2275] = c_Body_y[2274];
                    end else begin
                        n_Body_x[2275] = c_Body_x[c_Size-1];
                        n_Body_y[2275] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2276) begin
                        n_Body_x[2276] = c_Body_x[2275];
                        n_Body_y[2276] = c_Body_y[2275];
                    end else begin
                        n_Body_x[2276] = c_Body_x[c_Size-1];
                        n_Body_y[2276] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2277) begin
                        n_Body_x[2277] = c_Body_x[2276];
                        n_Body_y[2277] = c_Body_y[2276];
                    end else begin
                        n_Body_x[2277] = c_Body_x[c_Size-1];
                        n_Body_y[2277] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2278) begin
                        n_Body_x[2278] = c_Body_x[2277];
                        n_Body_y[2278] = c_Body_y[2277];
                    end else begin
                        n_Body_x[2278] = c_Body_x[c_Size-1];
                        n_Body_y[2278] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2279) begin
                        n_Body_x[2279] = c_Body_x[2278];
                        n_Body_y[2279] = c_Body_y[2278];
                    end else begin
                        n_Body_x[2279] = c_Body_x[c_Size-1];
                        n_Body_y[2279] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2280) begin
                        n_Body_x[2280] = c_Body_x[2279];
                        n_Body_y[2280] = c_Body_y[2279];
                    end else begin
                        n_Body_x[2280] = c_Body_x[c_Size-1];
                        n_Body_y[2280] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2281) begin
                        n_Body_x[2281] = c_Body_x[2280];
                        n_Body_y[2281] = c_Body_y[2280];
                    end else begin
                        n_Body_x[2281] = c_Body_x[c_Size-1];
                        n_Body_y[2281] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2282) begin
                        n_Body_x[2282] = c_Body_x[2281];
                        n_Body_y[2282] = c_Body_y[2281];
                    end else begin
                        n_Body_x[2282] = c_Body_x[c_Size-1];
                        n_Body_y[2282] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2283) begin
                        n_Body_x[2283] = c_Body_x[2282];
                        n_Body_y[2283] = c_Body_y[2282];
                    end else begin
                        n_Body_x[2283] = c_Body_x[c_Size-1];
                        n_Body_y[2283] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2284) begin
                        n_Body_x[2284] = c_Body_x[2283];
                        n_Body_y[2284] = c_Body_y[2283];
                    end else begin
                        n_Body_x[2284] = c_Body_x[c_Size-1];
                        n_Body_y[2284] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2285) begin
                        n_Body_x[2285] = c_Body_x[2284];
                        n_Body_y[2285] = c_Body_y[2284];
                    end else begin
                        n_Body_x[2285] = c_Body_x[c_Size-1];
                        n_Body_y[2285] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2286) begin
                        n_Body_x[2286] = c_Body_x[2285];
                        n_Body_y[2286] = c_Body_y[2285];
                    end else begin
                        n_Body_x[2286] = c_Body_x[c_Size-1];
                        n_Body_y[2286] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2287) begin
                        n_Body_x[2287] = c_Body_x[2286];
                        n_Body_y[2287] = c_Body_y[2286];
                    end else begin
                        n_Body_x[2287] = c_Body_x[c_Size-1];
                        n_Body_y[2287] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2288) begin
                        n_Body_x[2288] = c_Body_x[2287];
                        n_Body_y[2288] = c_Body_y[2287];
                    end else begin
                        n_Body_x[2288] = c_Body_x[c_Size-1];
                        n_Body_y[2288] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2289) begin
                        n_Body_x[2289] = c_Body_x[2288];
                        n_Body_y[2289] = c_Body_y[2288];
                    end else begin
                        n_Body_x[2289] = c_Body_x[c_Size-1];
                        n_Body_y[2289] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2290) begin
                        n_Body_x[2290] = c_Body_x[2289];
                        n_Body_y[2290] = c_Body_y[2289];
                    end else begin
                        n_Body_x[2290] = c_Body_x[c_Size-1];
                        n_Body_y[2290] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2291) begin
                        n_Body_x[2291] = c_Body_x[2290];
                        n_Body_y[2291] = c_Body_y[2290];
                    end else begin
                        n_Body_x[2291] = c_Body_x[c_Size-1];
                        n_Body_y[2291] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2292) begin
                        n_Body_x[2292] = c_Body_x[2291];
                        n_Body_y[2292] = c_Body_y[2291];
                    end else begin
                        n_Body_x[2292] = c_Body_x[c_Size-1];
                        n_Body_y[2292] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2293) begin
                        n_Body_x[2293] = c_Body_x[2292];
                        n_Body_y[2293] = c_Body_y[2292];
                    end else begin
                        n_Body_x[2293] = c_Body_x[c_Size-1];
                        n_Body_y[2293] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2294) begin
                        n_Body_x[2294] = c_Body_x[2293];
                        n_Body_y[2294] = c_Body_y[2293];
                    end else begin
                        n_Body_x[2294] = c_Body_x[c_Size-1];
                        n_Body_y[2294] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2295) begin
                        n_Body_x[2295] = c_Body_x[2294];
                        n_Body_y[2295] = c_Body_y[2294];
                    end else begin
                        n_Body_x[2295] = c_Body_x[c_Size-1];
                        n_Body_y[2295] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2296) begin
                        n_Body_x[2296] = c_Body_x[2295];
                        n_Body_y[2296] = c_Body_y[2295];
                    end else begin
                        n_Body_x[2296] = c_Body_x[c_Size-1];
                        n_Body_y[2296] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2297) begin
                        n_Body_x[2297] = c_Body_x[2296];
                        n_Body_y[2297] = c_Body_y[2296];
                    end else begin
                        n_Body_x[2297] = c_Body_x[c_Size-1];
                        n_Body_y[2297] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2298) begin
                        n_Body_x[2298] = c_Body_x[2297];
                        n_Body_y[2298] = c_Body_y[2297];
                    end else begin
                        n_Body_x[2298] = c_Body_x[c_Size-1];
                        n_Body_y[2298] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2299) begin
                        n_Body_x[2299] = c_Body_x[2298];
                        n_Body_y[2299] = c_Body_y[2298];
                    end else begin
                        n_Body_x[2299] = c_Body_x[c_Size-1];
                        n_Body_y[2299] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2300) begin
                        n_Body_x[2300] = c_Body_x[2299];
                        n_Body_y[2300] = c_Body_y[2299];
                    end else begin
                        n_Body_x[2300] = c_Body_x[c_Size-1];
                        n_Body_y[2300] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2301) begin
                        n_Body_x[2301] = c_Body_x[2300];
                        n_Body_y[2301] = c_Body_y[2300];
                    end else begin
                        n_Body_x[2301] = c_Body_x[c_Size-1];
                        n_Body_y[2301] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2302) begin
                        n_Body_x[2302] = c_Body_x[2301];
                        n_Body_y[2302] = c_Body_y[2301];
                    end else begin
                        n_Body_x[2302] = c_Body_x[c_Size-1];
                        n_Body_y[2302] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2303) begin
                        n_Body_x[2303] = c_Body_x[2302];
                        n_Body_y[2303] = c_Body_y[2302];
                    end else begin
                        n_Body_x[2303] = c_Body_x[c_Size-1];
                        n_Body_y[2303] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2304) begin
                        n_Body_x[2304] = c_Body_x[2303];
                        n_Body_y[2304] = c_Body_y[2303];
                    end else begin
                        n_Body_x[2304] = c_Body_x[c_Size-1];
                        n_Body_y[2304] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2305) begin
                        n_Body_x[2305] = c_Body_x[2304];
                        n_Body_y[2305] = c_Body_y[2304];
                    end else begin
                        n_Body_x[2305] = c_Body_x[c_Size-1];
                        n_Body_y[2305] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2306) begin
                        n_Body_x[2306] = c_Body_x[2305];
                        n_Body_y[2306] = c_Body_y[2305];
                    end else begin
                        n_Body_x[2306] = c_Body_x[c_Size-1];
                        n_Body_y[2306] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2307) begin
                        n_Body_x[2307] = c_Body_x[2306];
                        n_Body_y[2307] = c_Body_y[2306];
                    end else begin
                        n_Body_x[2307] = c_Body_x[c_Size-1];
                        n_Body_y[2307] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2308) begin
                        n_Body_x[2308] = c_Body_x[2307];
                        n_Body_y[2308] = c_Body_y[2307];
                    end else begin
                        n_Body_x[2308] = c_Body_x[c_Size-1];
                        n_Body_y[2308] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2309) begin
                        n_Body_x[2309] = c_Body_x[2308];
                        n_Body_y[2309] = c_Body_y[2308];
                    end else begin
                        n_Body_x[2309] = c_Body_x[c_Size-1];
                        n_Body_y[2309] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2310) begin
                        n_Body_x[2310] = c_Body_x[2309];
                        n_Body_y[2310] = c_Body_y[2309];
                    end else begin
                        n_Body_x[2310] = c_Body_x[c_Size-1];
                        n_Body_y[2310] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2311) begin
                        n_Body_x[2311] = c_Body_x[2310];
                        n_Body_y[2311] = c_Body_y[2310];
                    end else begin
                        n_Body_x[2311] = c_Body_x[c_Size-1];
                        n_Body_y[2311] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2312) begin
                        n_Body_x[2312] = c_Body_x[2311];
                        n_Body_y[2312] = c_Body_y[2311];
                    end else begin
                        n_Body_x[2312] = c_Body_x[c_Size-1];
                        n_Body_y[2312] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2313) begin
                        n_Body_x[2313] = c_Body_x[2312];
                        n_Body_y[2313] = c_Body_y[2312];
                    end else begin
                        n_Body_x[2313] = c_Body_x[c_Size-1];
                        n_Body_y[2313] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2314) begin
                        n_Body_x[2314] = c_Body_x[2313];
                        n_Body_y[2314] = c_Body_y[2313];
                    end else begin
                        n_Body_x[2314] = c_Body_x[c_Size-1];
                        n_Body_y[2314] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2315) begin
                        n_Body_x[2315] = c_Body_x[2314];
                        n_Body_y[2315] = c_Body_y[2314];
                    end else begin
                        n_Body_x[2315] = c_Body_x[c_Size-1];
                        n_Body_y[2315] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2316) begin
                        n_Body_x[2316] = c_Body_x[2315];
                        n_Body_y[2316] = c_Body_y[2315];
                    end else begin
                        n_Body_x[2316] = c_Body_x[c_Size-1];
                        n_Body_y[2316] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2317) begin
                        n_Body_x[2317] = c_Body_x[2316];
                        n_Body_y[2317] = c_Body_y[2316];
                    end else begin
                        n_Body_x[2317] = c_Body_x[c_Size-1];
                        n_Body_y[2317] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2318) begin
                        n_Body_x[2318] = c_Body_x[2317];
                        n_Body_y[2318] = c_Body_y[2317];
                    end else begin
                        n_Body_x[2318] = c_Body_x[c_Size-1];
                        n_Body_y[2318] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2319) begin
                        n_Body_x[2319] = c_Body_x[2318];
                        n_Body_y[2319] = c_Body_y[2318];
                    end else begin
                        n_Body_x[2319] = c_Body_x[c_Size-1];
                        n_Body_y[2319] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2320) begin
                        n_Body_x[2320] = c_Body_x[2319];
                        n_Body_y[2320] = c_Body_y[2319];
                    end else begin
                        n_Body_x[2320] = c_Body_x[c_Size-1];
                        n_Body_y[2320] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2321) begin
                        n_Body_x[2321] = c_Body_x[2320];
                        n_Body_y[2321] = c_Body_y[2320];
                    end else begin
                        n_Body_x[2321] = c_Body_x[c_Size-1];
                        n_Body_y[2321] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2322) begin
                        n_Body_x[2322] = c_Body_x[2321];
                        n_Body_y[2322] = c_Body_y[2321];
                    end else begin
                        n_Body_x[2322] = c_Body_x[c_Size-1];
                        n_Body_y[2322] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2323) begin
                        n_Body_x[2323] = c_Body_x[2322];
                        n_Body_y[2323] = c_Body_y[2322];
                    end else begin
                        n_Body_x[2323] = c_Body_x[c_Size-1];
                        n_Body_y[2323] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2324) begin
                        n_Body_x[2324] = c_Body_x[2323];
                        n_Body_y[2324] = c_Body_y[2323];
                    end else begin
                        n_Body_x[2324] = c_Body_x[c_Size-1];
                        n_Body_y[2324] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2325) begin
                        n_Body_x[2325] = c_Body_x[2324];
                        n_Body_y[2325] = c_Body_y[2324];
                    end else begin
                        n_Body_x[2325] = c_Body_x[c_Size-1];
                        n_Body_y[2325] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2326) begin
                        n_Body_x[2326] = c_Body_x[2325];
                        n_Body_y[2326] = c_Body_y[2325];
                    end else begin
                        n_Body_x[2326] = c_Body_x[c_Size-1];
                        n_Body_y[2326] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2327) begin
                        n_Body_x[2327] = c_Body_x[2326];
                        n_Body_y[2327] = c_Body_y[2326];
                    end else begin
                        n_Body_x[2327] = c_Body_x[c_Size-1];
                        n_Body_y[2327] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2328) begin
                        n_Body_x[2328] = c_Body_x[2327];
                        n_Body_y[2328] = c_Body_y[2327];
                    end else begin
                        n_Body_x[2328] = c_Body_x[c_Size-1];
                        n_Body_y[2328] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2329) begin
                        n_Body_x[2329] = c_Body_x[2328];
                        n_Body_y[2329] = c_Body_y[2328];
                    end else begin
                        n_Body_x[2329] = c_Body_x[c_Size-1];
                        n_Body_y[2329] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2330) begin
                        n_Body_x[2330] = c_Body_x[2329];
                        n_Body_y[2330] = c_Body_y[2329];
                    end else begin
                        n_Body_x[2330] = c_Body_x[c_Size-1];
                        n_Body_y[2330] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2331) begin
                        n_Body_x[2331] = c_Body_x[2330];
                        n_Body_y[2331] = c_Body_y[2330];
                    end else begin
                        n_Body_x[2331] = c_Body_x[c_Size-1];
                        n_Body_y[2331] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2332) begin
                        n_Body_x[2332] = c_Body_x[2331];
                        n_Body_y[2332] = c_Body_y[2331];
                    end else begin
                        n_Body_x[2332] = c_Body_x[c_Size-1];
                        n_Body_y[2332] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2333) begin
                        n_Body_x[2333] = c_Body_x[2332];
                        n_Body_y[2333] = c_Body_y[2332];
                    end else begin
                        n_Body_x[2333] = c_Body_x[c_Size-1];
                        n_Body_y[2333] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2334) begin
                        n_Body_x[2334] = c_Body_x[2333];
                        n_Body_y[2334] = c_Body_y[2333];
                    end else begin
                        n_Body_x[2334] = c_Body_x[c_Size-1];
                        n_Body_y[2334] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2335) begin
                        n_Body_x[2335] = c_Body_x[2334];
                        n_Body_y[2335] = c_Body_y[2334];
                    end else begin
                        n_Body_x[2335] = c_Body_x[c_Size-1];
                        n_Body_y[2335] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2336) begin
                        n_Body_x[2336] = c_Body_x[2335];
                        n_Body_y[2336] = c_Body_y[2335];
                    end else begin
                        n_Body_x[2336] = c_Body_x[c_Size-1];
                        n_Body_y[2336] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2337) begin
                        n_Body_x[2337] = c_Body_x[2336];
                        n_Body_y[2337] = c_Body_y[2336];
                    end else begin
                        n_Body_x[2337] = c_Body_x[c_Size-1];
                        n_Body_y[2337] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2338) begin
                        n_Body_x[2338] = c_Body_x[2337];
                        n_Body_y[2338] = c_Body_y[2337];
                    end else begin
                        n_Body_x[2338] = c_Body_x[c_Size-1];
                        n_Body_y[2338] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2339) begin
                        n_Body_x[2339] = c_Body_x[2338];
                        n_Body_y[2339] = c_Body_y[2338];
                    end else begin
                        n_Body_x[2339] = c_Body_x[c_Size-1];
                        n_Body_y[2339] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2340) begin
                        n_Body_x[2340] = c_Body_x[2339];
                        n_Body_y[2340] = c_Body_y[2339];
                    end else begin
                        n_Body_x[2340] = c_Body_x[c_Size-1];
                        n_Body_y[2340] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2341) begin
                        n_Body_x[2341] = c_Body_x[2340];
                        n_Body_y[2341] = c_Body_y[2340];
                    end else begin
                        n_Body_x[2341] = c_Body_x[c_Size-1];
                        n_Body_y[2341] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2342) begin
                        n_Body_x[2342] = c_Body_x[2341];
                        n_Body_y[2342] = c_Body_y[2341];
                    end else begin
                        n_Body_x[2342] = c_Body_x[c_Size-1];
                        n_Body_y[2342] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2343) begin
                        n_Body_x[2343] = c_Body_x[2342];
                        n_Body_y[2343] = c_Body_y[2342];
                    end else begin
                        n_Body_x[2343] = c_Body_x[c_Size-1];
                        n_Body_y[2343] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2344) begin
                        n_Body_x[2344] = c_Body_x[2343];
                        n_Body_y[2344] = c_Body_y[2343];
                    end else begin
                        n_Body_x[2344] = c_Body_x[c_Size-1];
                        n_Body_y[2344] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2345) begin
                        n_Body_x[2345] = c_Body_x[2344];
                        n_Body_y[2345] = c_Body_y[2344];
                    end else begin
                        n_Body_x[2345] = c_Body_x[c_Size-1];
                        n_Body_y[2345] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2346) begin
                        n_Body_x[2346] = c_Body_x[2345];
                        n_Body_y[2346] = c_Body_y[2345];
                    end else begin
                        n_Body_x[2346] = c_Body_x[c_Size-1];
                        n_Body_y[2346] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2347) begin
                        n_Body_x[2347] = c_Body_x[2346];
                        n_Body_y[2347] = c_Body_y[2346];
                    end else begin
                        n_Body_x[2347] = c_Body_x[c_Size-1];
                        n_Body_y[2347] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2348) begin
                        n_Body_x[2348] = c_Body_x[2347];
                        n_Body_y[2348] = c_Body_y[2347];
                    end else begin
                        n_Body_x[2348] = c_Body_x[c_Size-1];
                        n_Body_y[2348] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2349) begin
                        n_Body_x[2349] = c_Body_x[2348];
                        n_Body_y[2349] = c_Body_y[2348];
                    end else begin
                        n_Body_x[2349] = c_Body_x[c_Size-1];
                        n_Body_y[2349] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2350) begin
                        n_Body_x[2350] = c_Body_x[2349];
                        n_Body_y[2350] = c_Body_y[2349];
                    end else begin
                        n_Body_x[2350] = c_Body_x[c_Size-1];
                        n_Body_y[2350] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2351) begin
                        n_Body_x[2351] = c_Body_x[2350];
                        n_Body_y[2351] = c_Body_y[2350];
                    end else begin
                        n_Body_x[2351] = c_Body_x[c_Size-1];
                        n_Body_y[2351] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2352) begin
                        n_Body_x[2352] = c_Body_x[2351];
                        n_Body_y[2352] = c_Body_y[2351];
                    end else begin
                        n_Body_x[2352] = c_Body_x[c_Size-1];
                        n_Body_y[2352] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2353) begin
                        n_Body_x[2353] = c_Body_x[2352];
                        n_Body_y[2353] = c_Body_y[2352];
                    end else begin
                        n_Body_x[2353] = c_Body_x[c_Size-1];
                        n_Body_y[2353] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2354) begin
                        n_Body_x[2354] = c_Body_x[2353];
                        n_Body_y[2354] = c_Body_y[2353];
                    end else begin
                        n_Body_x[2354] = c_Body_x[c_Size-1];
                        n_Body_y[2354] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2355) begin
                        n_Body_x[2355] = c_Body_x[2354];
                        n_Body_y[2355] = c_Body_y[2354];
                    end else begin
                        n_Body_x[2355] = c_Body_x[c_Size-1];
                        n_Body_y[2355] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2356) begin
                        n_Body_x[2356] = c_Body_x[2355];
                        n_Body_y[2356] = c_Body_y[2355];
                    end else begin
                        n_Body_x[2356] = c_Body_x[c_Size-1];
                        n_Body_y[2356] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2357) begin
                        n_Body_x[2357] = c_Body_x[2356];
                        n_Body_y[2357] = c_Body_y[2356];
                    end else begin
                        n_Body_x[2357] = c_Body_x[c_Size-1];
                        n_Body_y[2357] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2358) begin
                        n_Body_x[2358] = c_Body_x[2357];
                        n_Body_y[2358] = c_Body_y[2357];
                    end else begin
                        n_Body_x[2358] = c_Body_x[c_Size-1];
                        n_Body_y[2358] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2359) begin
                        n_Body_x[2359] = c_Body_x[2358];
                        n_Body_y[2359] = c_Body_y[2358];
                    end else begin
                        n_Body_x[2359] = c_Body_x[c_Size-1];
                        n_Body_y[2359] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2360) begin
                        n_Body_x[2360] = c_Body_x[2359];
                        n_Body_y[2360] = c_Body_y[2359];
                    end else begin
                        n_Body_x[2360] = c_Body_x[c_Size-1];
                        n_Body_y[2360] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2361) begin
                        n_Body_x[2361] = c_Body_x[2360];
                        n_Body_y[2361] = c_Body_y[2360];
                    end else begin
                        n_Body_x[2361] = c_Body_x[c_Size-1];
                        n_Body_y[2361] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2362) begin
                        n_Body_x[2362] = c_Body_x[2361];
                        n_Body_y[2362] = c_Body_y[2361];
                    end else begin
                        n_Body_x[2362] = c_Body_x[c_Size-1];
                        n_Body_y[2362] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2363) begin
                        n_Body_x[2363] = c_Body_x[2362];
                        n_Body_y[2363] = c_Body_y[2362];
                    end else begin
                        n_Body_x[2363] = c_Body_x[c_Size-1];
                        n_Body_y[2363] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2364) begin
                        n_Body_x[2364] = c_Body_x[2363];
                        n_Body_y[2364] = c_Body_y[2363];
                    end else begin
                        n_Body_x[2364] = c_Body_x[c_Size-1];
                        n_Body_y[2364] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2365) begin
                        n_Body_x[2365] = c_Body_x[2364];
                        n_Body_y[2365] = c_Body_y[2364];
                    end else begin
                        n_Body_x[2365] = c_Body_x[c_Size-1];
                        n_Body_y[2365] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2366) begin
                        n_Body_x[2366] = c_Body_x[2365];
                        n_Body_y[2366] = c_Body_y[2365];
                    end else begin
                        n_Body_x[2366] = c_Body_x[c_Size-1];
                        n_Body_y[2366] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2367) begin
                        n_Body_x[2367] = c_Body_x[2366];
                        n_Body_y[2367] = c_Body_y[2366];
                    end else begin
                        n_Body_x[2367] = c_Body_x[c_Size-1];
                        n_Body_y[2367] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2368) begin
                        n_Body_x[2368] = c_Body_x[2367];
                        n_Body_y[2368] = c_Body_y[2367];
                    end else begin
                        n_Body_x[2368] = c_Body_x[c_Size-1];
                        n_Body_y[2368] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2369) begin
                        n_Body_x[2369] = c_Body_x[2368];
                        n_Body_y[2369] = c_Body_y[2368];
                    end else begin
                        n_Body_x[2369] = c_Body_x[c_Size-1];
                        n_Body_y[2369] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2370) begin
                        n_Body_x[2370] = c_Body_x[2369];
                        n_Body_y[2370] = c_Body_y[2369];
                    end else begin
                        n_Body_x[2370] = c_Body_x[c_Size-1];
                        n_Body_y[2370] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2371) begin
                        n_Body_x[2371] = c_Body_x[2370];
                        n_Body_y[2371] = c_Body_y[2370];
                    end else begin
                        n_Body_x[2371] = c_Body_x[c_Size-1];
                        n_Body_y[2371] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2372) begin
                        n_Body_x[2372] = c_Body_x[2371];
                        n_Body_y[2372] = c_Body_y[2371];
                    end else begin
                        n_Body_x[2372] = c_Body_x[c_Size-1];
                        n_Body_y[2372] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2373) begin
                        n_Body_x[2373] = c_Body_x[2372];
                        n_Body_y[2373] = c_Body_y[2372];
                    end else begin
                        n_Body_x[2373] = c_Body_x[c_Size-1];
                        n_Body_y[2373] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2374) begin
                        n_Body_x[2374] = c_Body_x[2373];
                        n_Body_y[2374] = c_Body_y[2373];
                    end else begin
                        n_Body_x[2374] = c_Body_x[c_Size-1];
                        n_Body_y[2374] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2375) begin
                        n_Body_x[2375] = c_Body_x[2374];
                        n_Body_y[2375] = c_Body_y[2374];
                    end else begin
                        n_Body_x[2375] = c_Body_x[c_Size-1];
                        n_Body_y[2375] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2376) begin
                        n_Body_x[2376] = c_Body_x[2375];
                        n_Body_y[2376] = c_Body_y[2375];
                    end else begin
                        n_Body_x[2376] = c_Body_x[c_Size-1];
                        n_Body_y[2376] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2377) begin
                        n_Body_x[2377] = c_Body_x[2376];
                        n_Body_y[2377] = c_Body_y[2376];
                    end else begin
                        n_Body_x[2377] = c_Body_x[c_Size-1];
                        n_Body_y[2377] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2378) begin
                        n_Body_x[2378] = c_Body_x[2377];
                        n_Body_y[2378] = c_Body_y[2377];
                    end else begin
                        n_Body_x[2378] = c_Body_x[c_Size-1];
                        n_Body_y[2378] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2379) begin
                        n_Body_x[2379] = c_Body_x[2378];
                        n_Body_y[2379] = c_Body_y[2378];
                    end else begin
                        n_Body_x[2379] = c_Body_x[c_Size-1];
                        n_Body_y[2379] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2380) begin
                        n_Body_x[2380] = c_Body_x[2379];
                        n_Body_y[2380] = c_Body_y[2379];
                    end else begin
                        n_Body_x[2380] = c_Body_x[c_Size-1];
                        n_Body_y[2380] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2381) begin
                        n_Body_x[2381] = c_Body_x[2380];
                        n_Body_y[2381] = c_Body_y[2380];
                    end else begin
                        n_Body_x[2381] = c_Body_x[c_Size-1];
                        n_Body_y[2381] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2382) begin
                        n_Body_x[2382] = c_Body_x[2381];
                        n_Body_y[2382] = c_Body_y[2381];
                    end else begin
                        n_Body_x[2382] = c_Body_x[c_Size-1];
                        n_Body_y[2382] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2383) begin
                        n_Body_x[2383] = c_Body_x[2382];
                        n_Body_y[2383] = c_Body_y[2382];
                    end else begin
                        n_Body_x[2383] = c_Body_x[c_Size-1];
                        n_Body_y[2383] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2384) begin
                        n_Body_x[2384] = c_Body_x[2383];
                        n_Body_y[2384] = c_Body_y[2383];
                    end else begin
                        n_Body_x[2384] = c_Body_x[c_Size-1];
                        n_Body_y[2384] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2385) begin
                        n_Body_x[2385] = c_Body_x[2384];
                        n_Body_y[2385] = c_Body_y[2384];
                    end else begin
                        n_Body_x[2385] = c_Body_x[c_Size-1];
                        n_Body_y[2385] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2386) begin
                        n_Body_x[2386] = c_Body_x[2385];
                        n_Body_y[2386] = c_Body_y[2385];
                    end else begin
                        n_Body_x[2386] = c_Body_x[c_Size-1];
                        n_Body_y[2386] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2387) begin
                        n_Body_x[2387] = c_Body_x[2386];
                        n_Body_y[2387] = c_Body_y[2386];
                    end else begin
                        n_Body_x[2387] = c_Body_x[c_Size-1];
                        n_Body_y[2387] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2388) begin
                        n_Body_x[2388] = c_Body_x[2387];
                        n_Body_y[2388] = c_Body_y[2387];
                    end else begin
                        n_Body_x[2388] = c_Body_x[c_Size-1];
                        n_Body_y[2388] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2389) begin
                        n_Body_x[2389] = c_Body_x[2388];
                        n_Body_y[2389] = c_Body_y[2388];
                    end else begin
                        n_Body_x[2389] = c_Body_x[c_Size-1];
                        n_Body_y[2389] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2390) begin
                        n_Body_x[2390] = c_Body_x[2389];
                        n_Body_y[2390] = c_Body_y[2389];
                    end else begin
                        n_Body_x[2390] = c_Body_x[c_Size-1];
                        n_Body_y[2390] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2391) begin
                        n_Body_x[2391] = c_Body_x[2390];
                        n_Body_y[2391] = c_Body_y[2390];
                    end else begin
                        n_Body_x[2391] = c_Body_x[c_Size-1];
                        n_Body_y[2391] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2392) begin
                        n_Body_x[2392] = c_Body_x[2391];
                        n_Body_y[2392] = c_Body_y[2391];
                    end else begin
                        n_Body_x[2392] = c_Body_x[c_Size-1];
                        n_Body_y[2392] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2393) begin
                        n_Body_x[2393] = c_Body_x[2392];
                        n_Body_y[2393] = c_Body_y[2392];
                    end else begin
                        n_Body_x[2393] = c_Body_x[c_Size-1];
                        n_Body_y[2393] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2394) begin
                        n_Body_x[2394] = c_Body_x[2393];
                        n_Body_y[2394] = c_Body_y[2393];
                    end else begin
                        n_Body_x[2394] = c_Body_x[c_Size-1];
                        n_Body_y[2394] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2395) begin
                        n_Body_x[2395] = c_Body_x[2394];
                        n_Body_y[2395] = c_Body_y[2394];
                    end else begin
                        n_Body_x[2395] = c_Body_x[c_Size-1];
                        n_Body_y[2395] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2396) begin
                        n_Body_x[2396] = c_Body_x[2395];
                        n_Body_y[2396] = c_Body_y[2395];
                    end else begin
                        n_Body_x[2396] = c_Body_x[c_Size-1];
                        n_Body_y[2396] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2397) begin
                        n_Body_x[2397] = c_Body_x[2396];
                        n_Body_y[2397] = c_Body_y[2396];
                    end else begin
                        n_Body_x[2397] = c_Body_x[c_Size-1];
                        n_Body_y[2397] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2398) begin
                        n_Body_x[2398] = c_Body_x[2397];
                        n_Body_y[2398] = c_Body_y[2397];
                    end else begin
                        n_Body_x[2398] = c_Body_x[c_Size-1];
                        n_Body_y[2398] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2399) begin
                        n_Body_x[2399] = c_Body_x[2398];
                        n_Body_y[2399] = c_Body_y[2398];
                    end else begin
                        n_Body_x[2399] = c_Body_x[c_Size-1];
                        n_Body_y[2399] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2400) begin
                        n_Body_x[2400] = c_Body_x[2399];
                        n_Body_y[2400] = c_Body_y[2399];
                    end else begin
                        n_Body_x[2400] = c_Body_x[c_Size-1];
                        n_Body_y[2400] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2401) begin
                        n_Body_x[2401] = c_Body_x[2400];
                        n_Body_y[2401] = c_Body_y[2400];
                    end else begin
                        n_Body_x[2401] = c_Body_x[c_Size-1];
                        n_Body_y[2401] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2402) begin
                        n_Body_x[2402] = c_Body_x[2401];
                        n_Body_y[2402] = c_Body_y[2401];
                    end else begin
                        n_Body_x[2402] = c_Body_x[c_Size-1];
                        n_Body_y[2402] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2403) begin
                        n_Body_x[2403] = c_Body_x[2402];
                        n_Body_y[2403] = c_Body_y[2402];
                    end else begin
                        n_Body_x[2403] = c_Body_x[c_Size-1];
                        n_Body_y[2403] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2404) begin
                        n_Body_x[2404] = c_Body_x[2403];
                        n_Body_y[2404] = c_Body_y[2403];
                    end else begin
                        n_Body_x[2404] = c_Body_x[c_Size-1];
                        n_Body_y[2404] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2405) begin
                        n_Body_x[2405] = c_Body_x[2404];
                        n_Body_y[2405] = c_Body_y[2404];
                    end else begin
                        n_Body_x[2405] = c_Body_x[c_Size-1];
                        n_Body_y[2405] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2406) begin
                        n_Body_x[2406] = c_Body_x[2405];
                        n_Body_y[2406] = c_Body_y[2405];
                    end else begin
                        n_Body_x[2406] = c_Body_x[c_Size-1];
                        n_Body_y[2406] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2407) begin
                        n_Body_x[2407] = c_Body_x[2406];
                        n_Body_y[2407] = c_Body_y[2406];
                    end else begin
                        n_Body_x[2407] = c_Body_x[c_Size-1];
                        n_Body_y[2407] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2408) begin
                        n_Body_x[2408] = c_Body_x[2407];
                        n_Body_y[2408] = c_Body_y[2407];
                    end else begin
                        n_Body_x[2408] = c_Body_x[c_Size-1];
                        n_Body_y[2408] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2409) begin
                        n_Body_x[2409] = c_Body_x[2408];
                        n_Body_y[2409] = c_Body_y[2408];
                    end else begin
                        n_Body_x[2409] = c_Body_x[c_Size-1];
                        n_Body_y[2409] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2410) begin
                        n_Body_x[2410] = c_Body_x[2409];
                        n_Body_y[2410] = c_Body_y[2409];
                    end else begin
                        n_Body_x[2410] = c_Body_x[c_Size-1];
                        n_Body_y[2410] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2411) begin
                        n_Body_x[2411] = c_Body_x[2410];
                        n_Body_y[2411] = c_Body_y[2410];
                    end else begin
                        n_Body_x[2411] = c_Body_x[c_Size-1];
                        n_Body_y[2411] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2412) begin
                        n_Body_x[2412] = c_Body_x[2411];
                        n_Body_y[2412] = c_Body_y[2411];
                    end else begin
                        n_Body_x[2412] = c_Body_x[c_Size-1];
                        n_Body_y[2412] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2413) begin
                        n_Body_x[2413] = c_Body_x[2412];
                        n_Body_y[2413] = c_Body_y[2412];
                    end else begin
                        n_Body_x[2413] = c_Body_x[c_Size-1];
                        n_Body_y[2413] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2414) begin
                        n_Body_x[2414] = c_Body_x[2413];
                        n_Body_y[2414] = c_Body_y[2413];
                    end else begin
                        n_Body_x[2414] = c_Body_x[c_Size-1];
                        n_Body_y[2414] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2415) begin
                        n_Body_x[2415] = c_Body_x[2414];
                        n_Body_y[2415] = c_Body_y[2414];
                    end else begin
                        n_Body_x[2415] = c_Body_x[c_Size-1];
                        n_Body_y[2415] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2416) begin
                        n_Body_x[2416] = c_Body_x[2415];
                        n_Body_y[2416] = c_Body_y[2415];
                    end else begin
                        n_Body_x[2416] = c_Body_x[c_Size-1];
                        n_Body_y[2416] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2417) begin
                        n_Body_x[2417] = c_Body_x[2416];
                        n_Body_y[2417] = c_Body_y[2416];
                    end else begin
                        n_Body_x[2417] = c_Body_x[c_Size-1];
                        n_Body_y[2417] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2418) begin
                        n_Body_x[2418] = c_Body_x[2417];
                        n_Body_y[2418] = c_Body_y[2417];
                    end else begin
                        n_Body_x[2418] = c_Body_x[c_Size-1];
                        n_Body_y[2418] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2419) begin
                        n_Body_x[2419] = c_Body_x[2418];
                        n_Body_y[2419] = c_Body_y[2418];
                    end else begin
                        n_Body_x[2419] = c_Body_x[c_Size-1];
                        n_Body_y[2419] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2420) begin
                        n_Body_x[2420] = c_Body_x[2419];
                        n_Body_y[2420] = c_Body_y[2419];
                    end else begin
                        n_Body_x[2420] = c_Body_x[c_Size-1];
                        n_Body_y[2420] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2421) begin
                        n_Body_x[2421] = c_Body_x[2420];
                        n_Body_y[2421] = c_Body_y[2420];
                    end else begin
                        n_Body_x[2421] = c_Body_x[c_Size-1];
                        n_Body_y[2421] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2422) begin
                        n_Body_x[2422] = c_Body_x[2421];
                        n_Body_y[2422] = c_Body_y[2421];
                    end else begin
                        n_Body_x[2422] = c_Body_x[c_Size-1];
                        n_Body_y[2422] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2423) begin
                        n_Body_x[2423] = c_Body_x[2422];
                        n_Body_y[2423] = c_Body_y[2422];
                    end else begin
                        n_Body_x[2423] = c_Body_x[c_Size-1];
                        n_Body_y[2423] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2424) begin
                        n_Body_x[2424] = c_Body_x[2423];
                        n_Body_y[2424] = c_Body_y[2423];
                    end else begin
                        n_Body_x[2424] = c_Body_x[c_Size-1];
                        n_Body_y[2424] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2425) begin
                        n_Body_x[2425] = c_Body_x[2424];
                        n_Body_y[2425] = c_Body_y[2424];
                    end else begin
                        n_Body_x[2425] = c_Body_x[c_Size-1];
                        n_Body_y[2425] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2426) begin
                        n_Body_x[2426] = c_Body_x[2425];
                        n_Body_y[2426] = c_Body_y[2425];
                    end else begin
                        n_Body_x[2426] = c_Body_x[c_Size-1];
                        n_Body_y[2426] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2427) begin
                        n_Body_x[2427] = c_Body_x[2426];
                        n_Body_y[2427] = c_Body_y[2426];
                    end else begin
                        n_Body_x[2427] = c_Body_x[c_Size-1];
                        n_Body_y[2427] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2428) begin
                        n_Body_x[2428] = c_Body_x[2427];
                        n_Body_y[2428] = c_Body_y[2427];
                    end else begin
                        n_Body_x[2428] = c_Body_x[c_Size-1];
                        n_Body_y[2428] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2429) begin
                        n_Body_x[2429] = c_Body_x[2428];
                        n_Body_y[2429] = c_Body_y[2428];
                    end else begin
                        n_Body_x[2429] = c_Body_x[c_Size-1];
                        n_Body_y[2429] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2430) begin
                        n_Body_x[2430] = c_Body_x[2429];
                        n_Body_y[2430] = c_Body_y[2429];
                    end else begin
                        n_Body_x[2430] = c_Body_x[c_Size-1];
                        n_Body_y[2430] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2431) begin
                        n_Body_x[2431] = c_Body_x[2430];
                        n_Body_y[2431] = c_Body_y[2430];
                    end else begin
                        n_Body_x[2431] = c_Body_x[c_Size-1];
                        n_Body_y[2431] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2432) begin
                        n_Body_x[2432] = c_Body_x[2431];
                        n_Body_y[2432] = c_Body_y[2431];
                    end else begin
                        n_Body_x[2432] = c_Body_x[c_Size-1];
                        n_Body_y[2432] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2433) begin
                        n_Body_x[2433] = c_Body_x[2432];
                        n_Body_y[2433] = c_Body_y[2432];
                    end else begin
                        n_Body_x[2433] = c_Body_x[c_Size-1];
                        n_Body_y[2433] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2434) begin
                        n_Body_x[2434] = c_Body_x[2433];
                        n_Body_y[2434] = c_Body_y[2433];
                    end else begin
                        n_Body_x[2434] = c_Body_x[c_Size-1];
                        n_Body_y[2434] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2435) begin
                        n_Body_x[2435] = c_Body_x[2434];
                        n_Body_y[2435] = c_Body_y[2434];
                    end else begin
                        n_Body_x[2435] = c_Body_x[c_Size-1];
                        n_Body_y[2435] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2436) begin
                        n_Body_x[2436] = c_Body_x[2435];
                        n_Body_y[2436] = c_Body_y[2435];
                    end else begin
                        n_Body_x[2436] = c_Body_x[c_Size-1];
                        n_Body_y[2436] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2437) begin
                        n_Body_x[2437] = c_Body_x[2436];
                        n_Body_y[2437] = c_Body_y[2436];
                    end else begin
                        n_Body_x[2437] = c_Body_x[c_Size-1];
                        n_Body_y[2437] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2438) begin
                        n_Body_x[2438] = c_Body_x[2437];
                        n_Body_y[2438] = c_Body_y[2437];
                    end else begin
                        n_Body_x[2438] = c_Body_x[c_Size-1];
                        n_Body_y[2438] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2439) begin
                        n_Body_x[2439] = c_Body_x[2438];
                        n_Body_y[2439] = c_Body_y[2438];
                    end else begin
                        n_Body_x[2439] = c_Body_x[c_Size-1];
                        n_Body_y[2439] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2440) begin
                        n_Body_x[2440] = c_Body_x[2439];
                        n_Body_y[2440] = c_Body_y[2439];
                    end else begin
                        n_Body_x[2440] = c_Body_x[c_Size-1];
                        n_Body_y[2440] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2441) begin
                        n_Body_x[2441] = c_Body_x[2440];
                        n_Body_y[2441] = c_Body_y[2440];
                    end else begin
                        n_Body_x[2441] = c_Body_x[c_Size-1];
                        n_Body_y[2441] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2442) begin
                        n_Body_x[2442] = c_Body_x[2441];
                        n_Body_y[2442] = c_Body_y[2441];
                    end else begin
                        n_Body_x[2442] = c_Body_x[c_Size-1];
                        n_Body_y[2442] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2443) begin
                        n_Body_x[2443] = c_Body_x[2442];
                        n_Body_y[2443] = c_Body_y[2442];
                    end else begin
                        n_Body_x[2443] = c_Body_x[c_Size-1];
                        n_Body_y[2443] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2444) begin
                        n_Body_x[2444] = c_Body_x[2443];
                        n_Body_y[2444] = c_Body_y[2443];
                    end else begin
                        n_Body_x[2444] = c_Body_x[c_Size-1];
                        n_Body_y[2444] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2445) begin
                        n_Body_x[2445] = c_Body_x[2444];
                        n_Body_y[2445] = c_Body_y[2444];
                    end else begin
                        n_Body_x[2445] = c_Body_x[c_Size-1];
                        n_Body_y[2445] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2446) begin
                        n_Body_x[2446] = c_Body_x[2445];
                        n_Body_y[2446] = c_Body_y[2445];
                    end else begin
                        n_Body_x[2446] = c_Body_x[c_Size-1];
                        n_Body_y[2446] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2447) begin
                        n_Body_x[2447] = c_Body_x[2446];
                        n_Body_y[2447] = c_Body_y[2446];
                    end else begin
                        n_Body_x[2447] = c_Body_x[c_Size-1];
                        n_Body_y[2447] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2448) begin
                        n_Body_x[2448] = c_Body_x[2447];
                        n_Body_y[2448] = c_Body_y[2447];
                    end else begin
                        n_Body_x[2448] = c_Body_x[c_Size-1];
                        n_Body_y[2448] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2449) begin
                        n_Body_x[2449] = c_Body_x[2448];
                        n_Body_y[2449] = c_Body_y[2448];
                    end else begin
                        n_Body_x[2449] = c_Body_x[c_Size-1];
                        n_Body_y[2449] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2450) begin
                        n_Body_x[2450] = c_Body_x[2449];
                        n_Body_y[2450] = c_Body_y[2449];
                    end else begin
                        n_Body_x[2450] = c_Body_x[c_Size-1];
                        n_Body_y[2450] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2451) begin
                        n_Body_x[2451] = c_Body_x[2450];
                        n_Body_y[2451] = c_Body_y[2450];
                    end else begin
                        n_Body_x[2451] = c_Body_x[c_Size-1];
                        n_Body_y[2451] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2452) begin
                        n_Body_x[2452] = c_Body_x[2451];
                        n_Body_y[2452] = c_Body_y[2451];
                    end else begin
                        n_Body_x[2452] = c_Body_x[c_Size-1];
                        n_Body_y[2452] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2453) begin
                        n_Body_x[2453] = c_Body_x[2452];
                        n_Body_y[2453] = c_Body_y[2452];
                    end else begin
                        n_Body_x[2453] = c_Body_x[c_Size-1];
                        n_Body_y[2453] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2454) begin
                        n_Body_x[2454] = c_Body_x[2453];
                        n_Body_y[2454] = c_Body_y[2453];
                    end else begin
                        n_Body_x[2454] = c_Body_x[c_Size-1];
                        n_Body_y[2454] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2455) begin
                        n_Body_x[2455] = c_Body_x[2454];
                        n_Body_y[2455] = c_Body_y[2454];
                    end else begin
                        n_Body_x[2455] = c_Body_x[c_Size-1];
                        n_Body_y[2455] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2456) begin
                        n_Body_x[2456] = c_Body_x[2455];
                        n_Body_y[2456] = c_Body_y[2455];
                    end else begin
                        n_Body_x[2456] = c_Body_x[c_Size-1];
                        n_Body_y[2456] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2457) begin
                        n_Body_x[2457] = c_Body_x[2456];
                        n_Body_y[2457] = c_Body_y[2456];
                    end else begin
                        n_Body_x[2457] = c_Body_x[c_Size-1];
                        n_Body_y[2457] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2458) begin
                        n_Body_x[2458] = c_Body_x[2457];
                        n_Body_y[2458] = c_Body_y[2457];
                    end else begin
                        n_Body_x[2458] = c_Body_x[c_Size-1];
                        n_Body_y[2458] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2459) begin
                        n_Body_x[2459] = c_Body_x[2458];
                        n_Body_y[2459] = c_Body_y[2458];
                    end else begin
                        n_Body_x[2459] = c_Body_x[c_Size-1];
                        n_Body_y[2459] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2460) begin
                        n_Body_x[2460] = c_Body_x[2459];
                        n_Body_y[2460] = c_Body_y[2459];
                    end else begin
                        n_Body_x[2460] = c_Body_x[c_Size-1];
                        n_Body_y[2460] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2461) begin
                        n_Body_x[2461] = c_Body_x[2460];
                        n_Body_y[2461] = c_Body_y[2460];
                    end else begin
                        n_Body_x[2461] = c_Body_x[c_Size-1];
                        n_Body_y[2461] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2462) begin
                        n_Body_x[2462] = c_Body_x[2461];
                        n_Body_y[2462] = c_Body_y[2461];
                    end else begin
                        n_Body_x[2462] = c_Body_x[c_Size-1];
                        n_Body_y[2462] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2463) begin
                        n_Body_x[2463] = c_Body_x[2462];
                        n_Body_y[2463] = c_Body_y[2462];
                    end else begin
                        n_Body_x[2463] = c_Body_x[c_Size-1];
                        n_Body_y[2463] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2464) begin
                        n_Body_x[2464] = c_Body_x[2463];
                        n_Body_y[2464] = c_Body_y[2463];
                    end else begin
                        n_Body_x[2464] = c_Body_x[c_Size-1];
                        n_Body_y[2464] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2465) begin
                        n_Body_x[2465] = c_Body_x[2464];
                        n_Body_y[2465] = c_Body_y[2464];
                    end else begin
                        n_Body_x[2465] = c_Body_x[c_Size-1];
                        n_Body_y[2465] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2466) begin
                        n_Body_x[2466] = c_Body_x[2465];
                        n_Body_y[2466] = c_Body_y[2465];
                    end else begin
                        n_Body_x[2466] = c_Body_x[c_Size-1];
                        n_Body_y[2466] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2467) begin
                        n_Body_x[2467] = c_Body_x[2466];
                        n_Body_y[2467] = c_Body_y[2466];
                    end else begin
                        n_Body_x[2467] = c_Body_x[c_Size-1];
                        n_Body_y[2467] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2468) begin
                        n_Body_x[2468] = c_Body_x[2467];
                        n_Body_y[2468] = c_Body_y[2467];
                    end else begin
                        n_Body_x[2468] = c_Body_x[c_Size-1];
                        n_Body_y[2468] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2469) begin
                        n_Body_x[2469] = c_Body_x[2468];
                        n_Body_y[2469] = c_Body_y[2468];
                    end else begin
                        n_Body_x[2469] = c_Body_x[c_Size-1];
                        n_Body_y[2469] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2470) begin
                        n_Body_x[2470] = c_Body_x[2469];
                        n_Body_y[2470] = c_Body_y[2469];
                    end else begin
                        n_Body_x[2470] = c_Body_x[c_Size-1];
                        n_Body_y[2470] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2471) begin
                        n_Body_x[2471] = c_Body_x[2470];
                        n_Body_y[2471] = c_Body_y[2470];
                    end else begin
                        n_Body_x[2471] = c_Body_x[c_Size-1];
                        n_Body_y[2471] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2472) begin
                        n_Body_x[2472] = c_Body_x[2471];
                        n_Body_y[2472] = c_Body_y[2471];
                    end else begin
                        n_Body_x[2472] = c_Body_x[c_Size-1];
                        n_Body_y[2472] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2473) begin
                        n_Body_x[2473] = c_Body_x[2472];
                        n_Body_y[2473] = c_Body_y[2472];
                    end else begin
                        n_Body_x[2473] = c_Body_x[c_Size-1];
                        n_Body_y[2473] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2474) begin
                        n_Body_x[2474] = c_Body_x[2473];
                        n_Body_y[2474] = c_Body_y[2473];
                    end else begin
                        n_Body_x[2474] = c_Body_x[c_Size-1];
                        n_Body_y[2474] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2475) begin
                        n_Body_x[2475] = c_Body_x[2474];
                        n_Body_y[2475] = c_Body_y[2474];
                    end else begin
                        n_Body_x[2475] = c_Body_x[c_Size-1];
                        n_Body_y[2475] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2476) begin
                        n_Body_x[2476] = c_Body_x[2475];
                        n_Body_y[2476] = c_Body_y[2475];
                    end else begin
                        n_Body_x[2476] = c_Body_x[c_Size-1];
                        n_Body_y[2476] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2477) begin
                        n_Body_x[2477] = c_Body_x[2476];
                        n_Body_y[2477] = c_Body_y[2476];
                    end else begin
                        n_Body_x[2477] = c_Body_x[c_Size-1];
                        n_Body_y[2477] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2478) begin
                        n_Body_x[2478] = c_Body_x[2477];
                        n_Body_y[2478] = c_Body_y[2477];
                    end else begin
                        n_Body_x[2478] = c_Body_x[c_Size-1];
                        n_Body_y[2478] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2479) begin
                        n_Body_x[2479] = c_Body_x[2478];
                        n_Body_y[2479] = c_Body_y[2478];
                    end else begin
                        n_Body_x[2479] = c_Body_x[c_Size-1];
                        n_Body_y[2479] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2480) begin
                        n_Body_x[2480] = c_Body_x[2479];
                        n_Body_y[2480] = c_Body_y[2479];
                    end else begin
                        n_Body_x[2480] = c_Body_x[c_Size-1];
                        n_Body_y[2480] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2481) begin
                        n_Body_x[2481] = c_Body_x[2480];
                        n_Body_y[2481] = c_Body_y[2480];
                    end else begin
                        n_Body_x[2481] = c_Body_x[c_Size-1];
                        n_Body_y[2481] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2482) begin
                        n_Body_x[2482] = c_Body_x[2481];
                        n_Body_y[2482] = c_Body_y[2481];
                    end else begin
                        n_Body_x[2482] = c_Body_x[c_Size-1];
                        n_Body_y[2482] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2483) begin
                        n_Body_x[2483] = c_Body_x[2482];
                        n_Body_y[2483] = c_Body_y[2482];
                    end else begin
                        n_Body_x[2483] = c_Body_x[c_Size-1];
                        n_Body_y[2483] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2484) begin
                        n_Body_x[2484] = c_Body_x[2483];
                        n_Body_y[2484] = c_Body_y[2483];
                    end else begin
                        n_Body_x[2484] = c_Body_x[c_Size-1];
                        n_Body_y[2484] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2485) begin
                        n_Body_x[2485] = c_Body_x[2484];
                        n_Body_y[2485] = c_Body_y[2484];
                    end else begin
                        n_Body_x[2485] = c_Body_x[c_Size-1];
                        n_Body_y[2485] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2486) begin
                        n_Body_x[2486] = c_Body_x[2485];
                        n_Body_y[2486] = c_Body_y[2485];
                    end else begin
                        n_Body_x[2486] = c_Body_x[c_Size-1];
                        n_Body_y[2486] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2487) begin
                        n_Body_x[2487] = c_Body_x[2486];
                        n_Body_y[2487] = c_Body_y[2486];
                    end else begin
                        n_Body_x[2487] = c_Body_x[c_Size-1];
                        n_Body_y[2487] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2488) begin
                        n_Body_x[2488] = c_Body_x[2487];
                        n_Body_y[2488] = c_Body_y[2487];
                    end else begin
                        n_Body_x[2488] = c_Body_x[c_Size-1];
                        n_Body_y[2488] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2489) begin
                        n_Body_x[2489] = c_Body_x[2488];
                        n_Body_y[2489] = c_Body_y[2488];
                    end else begin
                        n_Body_x[2489] = c_Body_x[c_Size-1];
                        n_Body_y[2489] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2490) begin
                        n_Body_x[2490] = c_Body_x[2489];
                        n_Body_y[2490] = c_Body_y[2489];
                    end else begin
                        n_Body_x[2490] = c_Body_x[c_Size-1];
                        n_Body_y[2490] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2491) begin
                        n_Body_x[2491] = c_Body_x[2490];
                        n_Body_y[2491] = c_Body_y[2490];
                    end else begin
                        n_Body_x[2491] = c_Body_x[c_Size-1];
                        n_Body_y[2491] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2492) begin
                        n_Body_x[2492] = c_Body_x[2491];
                        n_Body_y[2492] = c_Body_y[2491];
                    end else begin
                        n_Body_x[2492] = c_Body_x[c_Size-1];
                        n_Body_y[2492] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2493) begin
                        n_Body_x[2493] = c_Body_x[2492];
                        n_Body_y[2493] = c_Body_y[2492];
                    end else begin
                        n_Body_x[2493] = c_Body_x[c_Size-1];
                        n_Body_y[2493] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2494) begin
                        n_Body_x[2494] = c_Body_x[2493];
                        n_Body_y[2494] = c_Body_y[2493];
                    end else begin
                        n_Body_x[2494] = c_Body_x[c_Size-1];
                        n_Body_y[2494] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2495) begin
                        n_Body_x[2495] = c_Body_x[2494];
                        n_Body_y[2495] = c_Body_y[2494];
                    end else begin
                        n_Body_x[2495] = c_Body_x[c_Size-1];
                        n_Body_y[2495] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2496) begin
                        n_Body_x[2496] = c_Body_x[2495];
                        n_Body_y[2496] = c_Body_y[2495];
                    end else begin
                        n_Body_x[2496] = c_Body_x[c_Size-1];
                        n_Body_y[2496] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2497) begin
                        n_Body_x[2497] = c_Body_x[2496];
                        n_Body_y[2497] = c_Body_y[2496];
                    end else begin
                        n_Body_x[2497] = c_Body_x[c_Size-1];
                        n_Body_y[2497] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2498) begin
                        n_Body_x[2498] = c_Body_x[2497];
                        n_Body_y[2498] = c_Body_y[2497];
                    end else begin
                        n_Body_x[2498] = c_Body_x[c_Size-1];
                        n_Body_y[2498] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2499) begin
                        n_Body_x[2499] = c_Body_x[2498];
                        n_Body_y[2499] = c_Body_y[2498];
                    end else begin
                        n_Body_x[2499] = c_Body_x[c_Size-1];
                        n_Body_y[2499] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2500) begin
                        n_Body_x[2500] = c_Body_x[2499];
                        n_Body_y[2500] = c_Body_y[2499];
                    end else begin
                        n_Body_x[2500] = c_Body_x[c_Size-1];
                        n_Body_y[2500] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2501) begin
                        n_Body_x[2501] = c_Body_x[2500];
                        n_Body_y[2501] = c_Body_y[2500];
                    end else begin
                        n_Body_x[2501] = c_Body_x[c_Size-1];
                        n_Body_y[2501] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2502) begin
                        n_Body_x[2502] = c_Body_x[2501];
                        n_Body_y[2502] = c_Body_y[2501];
                    end else begin
                        n_Body_x[2502] = c_Body_x[c_Size-1];
                        n_Body_y[2502] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2503) begin
                        n_Body_x[2503] = c_Body_x[2502];
                        n_Body_y[2503] = c_Body_y[2502];
                    end else begin
                        n_Body_x[2503] = c_Body_x[c_Size-1];
                        n_Body_y[2503] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2504) begin
                        n_Body_x[2504] = c_Body_x[2503];
                        n_Body_y[2504] = c_Body_y[2503];
                    end else begin
                        n_Body_x[2504] = c_Body_x[c_Size-1];
                        n_Body_y[2504] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2505) begin
                        n_Body_x[2505] = c_Body_x[2504];
                        n_Body_y[2505] = c_Body_y[2504];
                    end else begin
                        n_Body_x[2505] = c_Body_x[c_Size-1];
                        n_Body_y[2505] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2506) begin
                        n_Body_x[2506] = c_Body_x[2505];
                        n_Body_y[2506] = c_Body_y[2505];
                    end else begin
                        n_Body_x[2506] = c_Body_x[c_Size-1];
                        n_Body_y[2506] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2507) begin
                        n_Body_x[2507] = c_Body_x[2506];
                        n_Body_y[2507] = c_Body_y[2506];
                    end else begin
                        n_Body_x[2507] = c_Body_x[c_Size-1];
                        n_Body_y[2507] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2508) begin
                        n_Body_x[2508] = c_Body_x[2507];
                        n_Body_y[2508] = c_Body_y[2507];
                    end else begin
                        n_Body_x[2508] = c_Body_x[c_Size-1];
                        n_Body_y[2508] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2509) begin
                        n_Body_x[2509] = c_Body_x[2508];
                        n_Body_y[2509] = c_Body_y[2508];
                    end else begin
                        n_Body_x[2509] = c_Body_x[c_Size-1];
                        n_Body_y[2509] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2510) begin
                        n_Body_x[2510] = c_Body_x[2509];
                        n_Body_y[2510] = c_Body_y[2509];
                    end else begin
                        n_Body_x[2510] = c_Body_x[c_Size-1];
                        n_Body_y[2510] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2511) begin
                        n_Body_x[2511] = c_Body_x[2510];
                        n_Body_y[2511] = c_Body_y[2510];
                    end else begin
                        n_Body_x[2511] = c_Body_x[c_Size-1];
                        n_Body_y[2511] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2512) begin
                        n_Body_x[2512] = c_Body_x[2511];
                        n_Body_y[2512] = c_Body_y[2511];
                    end else begin
                        n_Body_x[2512] = c_Body_x[c_Size-1];
                        n_Body_y[2512] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2513) begin
                        n_Body_x[2513] = c_Body_x[2512];
                        n_Body_y[2513] = c_Body_y[2512];
                    end else begin
                        n_Body_x[2513] = c_Body_x[c_Size-1];
                        n_Body_y[2513] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2514) begin
                        n_Body_x[2514] = c_Body_x[2513];
                        n_Body_y[2514] = c_Body_y[2513];
                    end else begin
                        n_Body_x[2514] = c_Body_x[c_Size-1];
                        n_Body_y[2514] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2515) begin
                        n_Body_x[2515] = c_Body_x[2514];
                        n_Body_y[2515] = c_Body_y[2514];
                    end else begin
                        n_Body_x[2515] = c_Body_x[c_Size-1];
                        n_Body_y[2515] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2516) begin
                        n_Body_x[2516] = c_Body_x[2515];
                        n_Body_y[2516] = c_Body_y[2515];
                    end else begin
                        n_Body_x[2516] = c_Body_x[c_Size-1];
                        n_Body_y[2516] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2517) begin
                        n_Body_x[2517] = c_Body_x[2516];
                        n_Body_y[2517] = c_Body_y[2516];
                    end else begin
                        n_Body_x[2517] = c_Body_x[c_Size-1];
                        n_Body_y[2517] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2518) begin
                        n_Body_x[2518] = c_Body_x[2517];
                        n_Body_y[2518] = c_Body_y[2517];
                    end else begin
                        n_Body_x[2518] = c_Body_x[c_Size-1];
                        n_Body_y[2518] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2519) begin
                        n_Body_x[2519] = c_Body_x[2518];
                        n_Body_y[2519] = c_Body_y[2518];
                    end else begin
                        n_Body_x[2519] = c_Body_x[c_Size-1];
                        n_Body_y[2519] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2520) begin
                        n_Body_x[2520] = c_Body_x[2519];
                        n_Body_y[2520] = c_Body_y[2519];
                    end else begin
                        n_Body_x[2520] = c_Body_x[c_Size-1];
                        n_Body_y[2520] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2521) begin
                        n_Body_x[2521] = c_Body_x[2520];
                        n_Body_y[2521] = c_Body_y[2520];
                    end else begin
                        n_Body_x[2521] = c_Body_x[c_Size-1];
                        n_Body_y[2521] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2522) begin
                        n_Body_x[2522] = c_Body_x[2521];
                        n_Body_y[2522] = c_Body_y[2521];
                    end else begin
                        n_Body_x[2522] = c_Body_x[c_Size-1];
                        n_Body_y[2522] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2523) begin
                        n_Body_x[2523] = c_Body_x[2522];
                        n_Body_y[2523] = c_Body_y[2522];
                    end else begin
                        n_Body_x[2523] = c_Body_x[c_Size-1];
                        n_Body_y[2523] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2524) begin
                        n_Body_x[2524] = c_Body_x[2523];
                        n_Body_y[2524] = c_Body_y[2523];
                    end else begin
                        n_Body_x[2524] = c_Body_x[c_Size-1];
                        n_Body_y[2524] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2525) begin
                        n_Body_x[2525] = c_Body_x[2524];
                        n_Body_y[2525] = c_Body_y[2524];
                    end else begin
                        n_Body_x[2525] = c_Body_x[c_Size-1];
                        n_Body_y[2525] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2526) begin
                        n_Body_x[2526] = c_Body_x[2525];
                        n_Body_y[2526] = c_Body_y[2525];
                    end else begin
                        n_Body_x[2526] = c_Body_x[c_Size-1];
                        n_Body_y[2526] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2527) begin
                        n_Body_x[2527] = c_Body_x[2526];
                        n_Body_y[2527] = c_Body_y[2526];
                    end else begin
                        n_Body_x[2527] = c_Body_x[c_Size-1];
                        n_Body_y[2527] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2528) begin
                        n_Body_x[2528] = c_Body_x[2527];
                        n_Body_y[2528] = c_Body_y[2527];
                    end else begin
                        n_Body_x[2528] = c_Body_x[c_Size-1];
                        n_Body_y[2528] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2529) begin
                        n_Body_x[2529] = c_Body_x[2528];
                        n_Body_y[2529] = c_Body_y[2528];
                    end else begin
                        n_Body_x[2529] = c_Body_x[c_Size-1];
                        n_Body_y[2529] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2530) begin
                        n_Body_x[2530] = c_Body_x[2529];
                        n_Body_y[2530] = c_Body_y[2529];
                    end else begin
                        n_Body_x[2530] = c_Body_x[c_Size-1];
                        n_Body_y[2530] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2531) begin
                        n_Body_x[2531] = c_Body_x[2530];
                        n_Body_y[2531] = c_Body_y[2530];
                    end else begin
                        n_Body_x[2531] = c_Body_x[c_Size-1];
                        n_Body_y[2531] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2532) begin
                        n_Body_x[2532] = c_Body_x[2531];
                        n_Body_y[2532] = c_Body_y[2531];
                    end else begin
                        n_Body_x[2532] = c_Body_x[c_Size-1];
                        n_Body_y[2532] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2533) begin
                        n_Body_x[2533] = c_Body_x[2532];
                        n_Body_y[2533] = c_Body_y[2532];
                    end else begin
                        n_Body_x[2533] = c_Body_x[c_Size-1];
                        n_Body_y[2533] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2534) begin
                        n_Body_x[2534] = c_Body_x[2533];
                        n_Body_y[2534] = c_Body_y[2533];
                    end else begin
                        n_Body_x[2534] = c_Body_x[c_Size-1];
                        n_Body_y[2534] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2535) begin
                        n_Body_x[2535] = c_Body_x[2534];
                        n_Body_y[2535] = c_Body_y[2534];
                    end else begin
                        n_Body_x[2535] = c_Body_x[c_Size-1];
                        n_Body_y[2535] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2536) begin
                        n_Body_x[2536] = c_Body_x[2535];
                        n_Body_y[2536] = c_Body_y[2535];
                    end else begin
                        n_Body_x[2536] = c_Body_x[c_Size-1];
                        n_Body_y[2536] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2537) begin
                        n_Body_x[2537] = c_Body_x[2536];
                        n_Body_y[2537] = c_Body_y[2536];
                    end else begin
                        n_Body_x[2537] = c_Body_x[c_Size-1];
                        n_Body_y[2537] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2538) begin
                        n_Body_x[2538] = c_Body_x[2537];
                        n_Body_y[2538] = c_Body_y[2537];
                    end else begin
                        n_Body_x[2538] = c_Body_x[c_Size-1];
                        n_Body_y[2538] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2539) begin
                        n_Body_x[2539] = c_Body_x[2538];
                        n_Body_y[2539] = c_Body_y[2538];
                    end else begin
                        n_Body_x[2539] = c_Body_x[c_Size-1];
                        n_Body_y[2539] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2540) begin
                        n_Body_x[2540] = c_Body_x[2539];
                        n_Body_y[2540] = c_Body_y[2539];
                    end else begin
                        n_Body_x[2540] = c_Body_x[c_Size-1];
                        n_Body_y[2540] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2541) begin
                        n_Body_x[2541] = c_Body_x[2540];
                        n_Body_y[2541] = c_Body_y[2540];
                    end else begin
                        n_Body_x[2541] = c_Body_x[c_Size-1];
                        n_Body_y[2541] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2542) begin
                        n_Body_x[2542] = c_Body_x[2541];
                        n_Body_y[2542] = c_Body_y[2541];
                    end else begin
                        n_Body_x[2542] = c_Body_x[c_Size-1];
                        n_Body_y[2542] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2543) begin
                        n_Body_x[2543] = c_Body_x[2542];
                        n_Body_y[2543] = c_Body_y[2542];
                    end else begin
                        n_Body_x[2543] = c_Body_x[c_Size-1];
                        n_Body_y[2543] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2544) begin
                        n_Body_x[2544] = c_Body_x[2543];
                        n_Body_y[2544] = c_Body_y[2543];
                    end else begin
                        n_Body_x[2544] = c_Body_x[c_Size-1];
                        n_Body_y[2544] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2545) begin
                        n_Body_x[2545] = c_Body_x[2544];
                        n_Body_y[2545] = c_Body_y[2544];
                    end else begin
                        n_Body_x[2545] = c_Body_x[c_Size-1];
                        n_Body_y[2545] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2546) begin
                        n_Body_x[2546] = c_Body_x[2545];
                        n_Body_y[2546] = c_Body_y[2545];
                    end else begin
                        n_Body_x[2546] = c_Body_x[c_Size-1];
                        n_Body_y[2546] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2547) begin
                        n_Body_x[2547] = c_Body_x[2546];
                        n_Body_y[2547] = c_Body_y[2546];
                    end else begin
                        n_Body_x[2547] = c_Body_x[c_Size-1];
                        n_Body_y[2547] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2548) begin
                        n_Body_x[2548] = c_Body_x[2547];
                        n_Body_y[2548] = c_Body_y[2547];
                    end else begin
                        n_Body_x[2548] = c_Body_x[c_Size-1];
                        n_Body_y[2548] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2549) begin
                        n_Body_x[2549] = c_Body_x[2548];
                        n_Body_y[2549] = c_Body_y[2548];
                    end else begin
                        n_Body_x[2549] = c_Body_x[c_Size-1];
                        n_Body_y[2549] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2550) begin
                        n_Body_x[2550] = c_Body_x[2549];
                        n_Body_y[2550] = c_Body_y[2549];
                    end else begin
                        n_Body_x[2550] = c_Body_x[c_Size-1];
                        n_Body_y[2550] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2551) begin
                        n_Body_x[2551] = c_Body_x[2550];
                        n_Body_y[2551] = c_Body_y[2550];
                    end else begin
                        n_Body_x[2551] = c_Body_x[c_Size-1];
                        n_Body_y[2551] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2552) begin
                        n_Body_x[2552] = c_Body_x[2551];
                        n_Body_y[2552] = c_Body_y[2551];
                    end else begin
                        n_Body_x[2552] = c_Body_x[c_Size-1];
                        n_Body_y[2552] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2553) begin
                        n_Body_x[2553] = c_Body_x[2552];
                        n_Body_y[2553] = c_Body_y[2552];
                    end else begin
                        n_Body_x[2553] = c_Body_x[c_Size-1];
                        n_Body_y[2553] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2554) begin
                        n_Body_x[2554] = c_Body_x[2553];
                        n_Body_y[2554] = c_Body_y[2553];
                    end else begin
                        n_Body_x[2554] = c_Body_x[c_Size-1];
                        n_Body_y[2554] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2555) begin
                        n_Body_x[2555] = c_Body_x[2554];
                        n_Body_y[2555] = c_Body_y[2554];
                    end else begin
                        n_Body_x[2555] = c_Body_x[c_Size-1];
                        n_Body_y[2555] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2556) begin
                        n_Body_x[2556] = c_Body_x[2555];
                        n_Body_y[2556] = c_Body_y[2555];
                    end else begin
                        n_Body_x[2556] = c_Body_x[c_Size-1];
                        n_Body_y[2556] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2557) begin
                        n_Body_x[2557] = c_Body_x[2556];
                        n_Body_y[2557] = c_Body_y[2556];
                    end else begin
                        n_Body_x[2557] = c_Body_x[c_Size-1];
                        n_Body_y[2557] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2558) begin
                        n_Body_x[2558] = c_Body_x[2557];
                        n_Body_y[2558] = c_Body_y[2557];
                    end else begin
                        n_Body_x[2558] = c_Body_x[c_Size-1];
                        n_Body_y[2558] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2559) begin
                        n_Body_x[2559] = c_Body_x[2558];
                        n_Body_y[2559] = c_Body_y[2558];
                    end else begin
                        n_Body_x[2559] = c_Body_x[c_Size-1];
                        n_Body_y[2559] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2560) begin
                        n_Body_x[2560] = c_Body_x[2559];
                        n_Body_y[2560] = c_Body_y[2559];
                    end else begin
                        n_Body_x[2560] = c_Body_x[c_Size-1];
                        n_Body_y[2560] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2561) begin
                        n_Body_x[2561] = c_Body_x[2560];
                        n_Body_y[2561] = c_Body_y[2560];
                    end else begin
                        n_Body_x[2561] = c_Body_x[c_Size-1];
                        n_Body_y[2561] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2562) begin
                        n_Body_x[2562] = c_Body_x[2561];
                        n_Body_y[2562] = c_Body_y[2561];
                    end else begin
                        n_Body_x[2562] = c_Body_x[c_Size-1];
                        n_Body_y[2562] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2563) begin
                        n_Body_x[2563] = c_Body_x[2562];
                        n_Body_y[2563] = c_Body_y[2562];
                    end else begin
                        n_Body_x[2563] = c_Body_x[c_Size-1];
                        n_Body_y[2563] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2564) begin
                        n_Body_x[2564] = c_Body_x[2563];
                        n_Body_y[2564] = c_Body_y[2563];
                    end else begin
                        n_Body_x[2564] = c_Body_x[c_Size-1];
                        n_Body_y[2564] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2565) begin
                        n_Body_x[2565] = c_Body_x[2564];
                        n_Body_y[2565] = c_Body_y[2564];
                    end else begin
                        n_Body_x[2565] = c_Body_x[c_Size-1];
                        n_Body_y[2565] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2566) begin
                        n_Body_x[2566] = c_Body_x[2565];
                        n_Body_y[2566] = c_Body_y[2565];
                    end else begin
                        n_Body_x[2566] = c_Body_x[c_Size-1];
                        n_Body_y[2566] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2567) begin
                        n_Body_x[2567] = c_Body_x[2566];
                        n_Body_y[2567] = c_Body_y[2566];
                    end else begin
                        n_Body_x[2567] = c_Body_x[c_Size-1];
                        n_Body_y[2567] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2568) begin
                        n_Body_x[2568] = c_Body_x[2567];
                        n_Body_y[2568] = c_Body_y[2567];
                    end else begin
                        n_Body_x[2568] = c_Body_x[c_Size-1];
                        n_Body_y[2568] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2569) begin
                        n_Body_x[2569] = c_Body_x[2568];
                        n_Body_y[2569] = c_Body_y[2568];
                    end else begin
                        n_Body_x[2569] = c_Body_x[c_Size-1];
                        n_Body_y[2569] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2570) begin
                        n_Body_x[2570] = c_Body_x[2569];
                        n_Body_y[2570] = c_Body_y[2569];
                    end else begin
                        n_Body_x[2570] = c_Body_x[c_Size-1];
                        n_Body_y[2570] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2571) begin
                        n_Body_x[2571] = c_Body_x[2570];
                        n_Body_y[2571] = c_Body_y[2570];
                    end else begin
                        n_Body_x[2571] = c_Body_x[c_Size-1];
                        n_Body_y[2571] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2572) begin
                        n_Body_x[2572] = c_Body_x[2571];
                        n_Body_y[2572] = c_Body_y[2571];
                    end else begin
                        n_Body_x[2572] = c_Body_x[c_Size-1];
                        n_Body_y[2572] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2573) begin
                        n_Body_x[2573] = c_Body_x[2572];
                        n_Body_y[2573] = c_Body_y[2572];
                    end else begin
                        n_Body_x[2573] = c_Body_x[c_Size-1];
                        n_Body_y[2573] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2574) begin
                        n_Body_x[2574] = c_Body_x[2573];
                        n_Body_y[2574] = c_Body_y[2573];
                    end else begin
                        n_Body_x[2574] = c_Body_x[c_Size-1];
                        n_Body_y[2574] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2575) begin
                        n_Body_x[2575] = c_Body_x[2574];
                        n_Body_y[2575] = c_Body_y[2574];
                    end else begin
                        n_Body_x[2575] = c_Body_x[c_Size-1];
                        n_Body_y[2575] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2576) begin
                        n_Body_x[2576] = c_Body_x[2575];
                        n_Body_y[2576] = c_Body_y[2575];
                    end else begin
                        n_Body_x[2576] = c_Body_x[c_Size-1];
                        n_Body_y[2576] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2577) begin
                        n_Body_x[2577] = c_Body_x[2576];
                        n_Body_y[2577] = c_Body_y[2576];
                    end else begin
                        n_Body_x[2577] = c_Body_x[c_Size-1];
                        n_Body_y[2577] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2578) begin
                        n_Body_x[2578] = c_Body_x[2577];
                        n_Body_y[2578] = c_Body_y[2577];
                    end else begin
                        n_Body_x[2578] = c_Body_x[c_Size-1];
                        n_Body_y[2578] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2579) begin
                        n_Body_x[2579] = c_Body_x[2578];
                        n_Body_y[2579] = c_Body_y[2578];
                    end else begin
                        n_Body_x[2579] = c_Body_x[c_Size-1];
                        n_Body_y[2579] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2580) begin
                        n_Body_x[2580] = c_Body_x[2579];
                        n_Body_y[2580] = c_Body_y[2579];
                    end else begin
                        n_Body_x[2580] = c_Body_x[c_Size-1];
                        n_Body_y[2580] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2581) begin
                        n_Body_x[2581] = c_Body_x[2580];
                        n_Body_y[2581] = c_Body_y[2580];
                    end else begin
                        n_Body_x[2581] = c_Body_x[c_Size-1];
                        n_Body_y[2581] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2582) begin
                        n_Body_x[2582] = c_Body_x[2581];
                        n_Body_y[2582] = c_Body_y[2581];
                    end else begin
                        n_Body_x[2582] = c_Body_x[c_Size-1];
                        n_Body_y[2582] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2583) begin
                        n_Body_x[2583] = c_Body_x[2582];
                        n_Body_y[2583] = c_Body_y[2582];
                    end else begin
                        n_Body_x[2583] = c_Body_x[c_Size-1];
                        n_Body_y[2583] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2584) begin
                        n_Body_x[2584] = c_Body_x[2583];
                        n_Body_y[2584] = c_Body_y[2583];
                    end else begin
                        n_Body_x[2584] = c_Body_x[c_Size-1];
                        n_Body_y[2584] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2585) begin
                        n_Body_x[2585] = c_Body_x[2584];
                        n_Body_y[2585] = c_Body_y[2584];
                    end else begin
                        n_Body_x[2585] = c_Body_x[c_Size-1];
                        n_Body_y[2585] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2586) begin
                        n_Body_x[2586] = c_Body_x[2585];
                        n_Body_y[2586] = c_Body_y[2585];
                    end else begin
                        n_Body_x[2586] = c_Body_x[c_Size-1];
                        n_Body_y[2586] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2587) begin
                        n_Body_x[2587] = c_Body_x[2586];
                        n_Body_y[2587] = c_Body_y[2586];
                    end else begin
                        n_Body_x[2587] = c_Body_x[c_Size-1];
                        n_Body_y[2587] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2588) begin
                        n_Body_x[2588] = c_Body_x[2587];
                        n_Body_y[2588] = c_Body_y[2587];
                    end else begin
                        n_Body_x[2588] = c_Body_x[c_Size-1];
                        n_Body_y[2588] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2589) begin
                        n_Body_x[2589] = c_Body_x[2588];
                        n_Body_y[2589] = c_Body_y[2588];
                    end else begin
                        n_Body_x[2589] = c_Body_x[c_Size-1];
                        n_Body_y[2589] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2590) begin
                        n_Body_x[2590] = c_Body_x[2589];
                        n_Body_y[2590] = c_Body_y[2589];
                    end else begin
                        n_Body_x[2590] = c_Body_x[c_Size-1];
                        n_Body_y[2590] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2591) begin
                        n_Body_x[2591] = c_Body_x[2590];
                        n_Body_y[2591] = c_Body_y[2590];
                    end else begin
                        n_Body_x[2591] = c_Body_x[c_Size-1];
                        n_Body_y[2591] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2592) begin
                        n_Body_x[2592] = c_Body_x[2591];
                        n_Body_y[2592] = c_Body_y[2591];
                    end else begin
                        n_Body_x[2592] = c_Body_x[c_Size-1];
                        n_Body_y[2592] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2593) begin
                        n_Body_x[2593] = c_Body_x[2592];
                        n_Body_y[2593] = c_Body_y[2592];
                    end else begin
                        n_Body_x[2593] = c_Body_x[c_Size-1];
                        n_Body_y[2593] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2594) begin
                        n_Body_x[2594] = c_Body_x[2593];
                        n_Body_y[2594] = c_Body_y[2593];
                    end else begin
                        n_Body_x[2594] = c_Body_x[c_Size-1];
                        n_Body_y[2594] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2595) begin
                        n_Body_x[2595] = c_Body_x[2594];
                        n_Body_y[2595] = c_Body_y[2594];
                    end else begin
                        n_Body_x[2595] = c_Body_x[c_Size-1];
                        n_Body_y[2595] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2596) begin
                        n_Body_x[2596] = c_Body_x[2595];
                        n_Body_y[2596] = c_Body_y[2595];
                    end else begin
                        n_Body_x[2596] = c_Body_x[c_Size-1];
                        n_Body_y[2596] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2597) begin
                        n_Body_x[2597] = c_Body_x[2596];
                        n_Body_y[2597] = c_Body_y[2596];
                    end else begin
                        n_Body_x[2597] = c_Body_x[c_Size-1];
                        n_Body_y[2597] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2598) begin
                        n_Body_x[2598] = c_Body_x[2597];
                        n_Body_y[2598] = c_Body_y[2597];
                    end else begin
                        n_Body_x[2598] = c_Body_x[c_Size-1];
                        n_Body_y[2598] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2599) begin
                        n_Body_x[2599] = c_Body_x[2598];
                        n_Body_y[2599] = c_Body_y[2598];
                    end else begin
                        n_Body_x[2599] = c_Body_x[c_Size-1];
                        n_Body_y[2599] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2600) begin
                        n_Body_x[2600] = c_Body_x[2599];
                        n_Body_y[2600] = c_Body_y[2599];
                    end else begin
                        n_Body_x[2600] = c_Body_x[c_Size-1];
                        n_Body_y[2600] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2601) begin
                        n_Body_x[2601] = c_Body_x[2600];
                        n_Body_y[2601] = c_Body_y[2600];
                    end else begin
                        n_Body_x[2601] = c_Body_x[c_Size-1];
                        n_Body_y[2601] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2602) begin
                        n_Body_x[2602] = c_Body_x[2601];
                        n_Body_y[2602] = c_Body_y[2601];
                    end else begin
                        n_Body_x[2602] = c_Body_x[c_Size-1];
                        n_Body_y[2602] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2603) begin
                        n_Body_x[2603] = c_Body_x[2602];
                        n_Body_y[2603] = c_Body_y[2602];
                    end else begin
                        n_Body_x[2603] = c_Body_x[c_Size-1];
                        n_Body_y[2603] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2604) begin
                        n_Body_x[2604] = c_Body_x[2603];
                        n_Body_y[2604] = c_Body_y[2603];
                    end else begin
                        n_Body_x[2604] = c_Body_x[c_Size-1];
                        n_Body_y[2604] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2605) begin
                        n_Body_x[2605] = c_Body_x[2604];
                        n_Body_y[2605] = c_Body_y[2604];
                    end else begin
                        n_Body_x[2605] = c_Body_x[c_Size-1];
                        n_Body_y[2605] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2606) begin
                        n_Body_x[2606] = c_Body_x[2605];
                        n_Body_y[2606] = c_Body_y[2605];
                    end else begin
                        n_Body_x[2606] = c_Body_x[c_Size-1];
                        n_Body_y[2606] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2607) begin
                        n_Body_x[2607] = c_Body_x[2606];
                        n_Body_y[2607] = c_Body_y[2606];
                    end else begin
                        n_Body_x[2607] = c_Body_x[c_Size-1];
                        n_Body_y[2607] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2608) begin
                        n_Body_x[2608] = c_Body_x[2607];
                        n_Body_y[2608] = c_Body_y[2607];
                    end else begin
                        n_Body_x[2608] = c_Body_x[c_Size-1];
                        n_Body_y[2608] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2609) begin
                        n_Body_x[2609] = c_Body_x[2608];
                        n_Body_y[2609] = c_Body_y[2608];
                    end else begin
                        n_Body_x[2609] = c_Body_x[c_Size-1];
                        n_Body_y[2609] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2610) begin
                        n_Body_x[2610] = c_Body_x[2609];
                        n_Body_y[2610] = c_Body_y[2609];
                    end else begin
                        n_Body_x[2610] = c_Body_x[c_Size-1];
                        n_Body_y[2610] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2611) begin
                        n_Body_x[2611] = c_Body_x[2610];
                        n_Body_y[2611] = c_Body_y[2610];
                    end else begin
                        n_Body_x[2611] = c_Body_x[c_Size-1];
                        n_Body_y[2611] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2612) begin
                        n_Body_x[2612] = c_Body_x[2611];
                        n_Body_y[2612] = c_Body_y[2611];
                    end else begin
                        n_Body_x[2612] = c_Body_x[c_Size-1];
                        n_Body_y[2612] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2613) begin
                        n_Body_x[2613] = c_Body_x[2612];
                        n_Body_y[2613] = c_Body_y[2612];
                    end else begin
                        n_Body_x[2613] = c_Body_x[c_Size-1];
                        n_Body_y[2613] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2614) begin
                        n_Body_x[2614] = c_Body_x[2613];
                        n_Body_y[2614] = c_Body_y[2613];
                    end else begin
                        n_Body_x[2614] = c_Body_x[c_Size-1];
                        n_Body_y[2614] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2615) begin
                        n_Body_x[2615] = c_Body_x[2614];
                        n_Body_y[2615] = c_Body_y[2614];
                    end else begin
                        n_Body_x[2615] = c_Body_x[c_Size-1];
                        n_Body_y[2615] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2616) begin
                        n_Body_x[2616] = c_Body_x[2615];
                        n_Body_y[2616] = c_Body_y[2615];
                    end else begin
                        n_Body_x[2616] = c_Body_x[c_Size-1];
                        n_Body_y[2616] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2617) begin
                        n_Body_x[2617] = c_Body_x[2616];
                        n_Body_y[2617] = c_Body_y[2616];
                    end else begin
                        n_Body_x[2617] = c_Body_x[c_Size-1];
                        n_Body_y[2617] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2618) begin
                        n_Body_x[2618] = c_Body_x[2617];
                        n_Body_y[2618] = c_Body_y[2617];
                    end else begin
                        n_Body_x[2618] = c_Body_x[c_Size-1];
                        n_Body_y[2618] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2619) begin
                        n_Body_x[2619] = c_Body_x[2618];
                        n_Body_y[2619] = c_Body_y[2618];
                    end else begin
                        n_Body_x[2619] = c_Body_x[c_Size-1];
                        n_Body_y[2619] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2620) begin
                        n_Body_x[2620] = c_Body_x[2619];
                        n_Body_y[2620] = c_Body_y[2619];
                    end else begin
                        n_Body_x[2620] = c_Body_x[c_Size-1];
                        n_Body_y[2620] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2621) begin
                        n_Body_x[2621] = c_Body_x[2620];
                        n_Body_y[2621] = c_Body_y[2620];
                    end else begin
                        n_Body_x[2621] = c_Body_x[c_Size-1];
                        n_Body_y[2621] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2622) begin
                        n_Body_x[2622] = c_Body_x[2621];
                        n_Body_y[2622] = c_Body_y[2621];
                    end else begin
                        n_Body_x[2622] = c_Body_x[c_Size-1];
                        n_Body_y[2622] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2623) begin
                        n_Body_x[2623] = c_Body_x[2622];
                        n_Body_y[2623] = c_Body_y[2622];
                    end else begin
                        n_Body_x[2623] = c_Body_x[c_Size-1];
                        n_Body_y[2623] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2624) begin
                        n_Body_x[2624] = c_Body_x[2623];
                        n_Body_y[2624] = c_Body_y[2623];
                    end else begin
                        n_Body_x[2624] = c_Body_x[c_Size-1];
                        n_Body_y[2624] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2625) begin
                        n_Body_x[2625] = c_Body_x[2624];
                        n_Body_y[2625] = c_Body_y[2624];
                    end else begin
                        n_Body_x[2625] = c_Body_x[c_Size-1];
                        n_Body_y[2625] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2626) begin
                        n_Body_x[2626] = c_Body_x[2625];
                        n_Body_y[2626] = c_Body_y[2625];
                    end else begin
                        n_Body_x[2626] = c_Body_x[c_Size-1];
                        n_Body_y[2626] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2627) begin
                        n_Body_x[2627] = c_Body_x[2626];
                        n_Body_y[2627] = c_Body_y[2626];
                    end else begin
                        n_Body_x[2627] = c_Body_x[c_Size-1];
                        n_Body_y[2627] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2628) begin
                        n_Body_x[2628] = c_Body_x[2627];
                        n_Body_y[2628] = c_Body_y[2627];
                    end else begin
                        n_Body_x[2628] = c_Body_x[c_Size-1];
                        n_Body_y[2628] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2629) begin
                        n_Body_x[2629] = c_Body_x[2628];
                        n_Body_y[2629] = c_Body_y[2628];
                    end else begin
                        n_Body_x[2629] = c_Body_x[c_Size-1];
                        n_Body_y[2629] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2630) begin
                        n_Body_x[2630] = c_Body_x[2629];
                        n_Body_y[2630] = c_Body_y[2629];
                    end else begin
                        n_Body_x[2630] = c_Body_x[c_Size-1];
                        n_Body_y[2630] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2631) begin
                        n_Body_x[2631] = c_Body_x[2630];
                        n_Body_y[2631] = c_Body_y[2630];
                    end else begin
                        n_Body_x[2631] = c_Body_x[c_Size-1];
                        n_Body_y[2631] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2632) begin
                        n_Body_x[2632] = c_Body_x[2631];
                        n_Body_y[2632] = c_Body_y[2631];
                    end else begin
                        n_Body_x[2632] = c_Body_x[c_Size-1];
                        n_Body_y[2632] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2633) begin
                        n_Body_x[2633] = c_Body_x[2632];
                        n_Body_y[2633] = c_Body_y[2632];
                    end else begin
                        n_Body_x[2633] = c_Body_x[c_Size-1];
                        n_Body_y[2633] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2634) begin
                        n_Body_x[2634] = c_Body_x[2633];
                        n_Body_y[2634] = c_Body_y[2633];
                    end else begin
                        n_Body_x[2634] = c_Body_x[c_Size-1];
                        n_Body_y[2634] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2635) begin
                        n_Body_x[2635] = c_Body_x[2634];
                        n_Body_y[2635] = c_Body_y[2634];
                    end else begin
                        n_Body_x[2635] = c_Body_x[c_Size-1];
                        n_Body_y[2635] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2636) begin
                        n_Body_x[2636] = c_Body_x[2635];
                        n_Body_y[2636] = c_Body_y[2635];
                    end else begin
                        n_Body_x[2636] = c_Body_x[c_Size-1];
                        n_Body_y[2636] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2637) begin
                        n_Body_x[2637] = c_Body_x[2636];
                        n_Body_y[2637] = c_Body_y[2636];
                    end else begin
                        n_Body_x[2637] = c_Body_x[c_Size-1];
                        n_Body_y[2637] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2638) begin
                        n_Body_x[2638] = c_Body_x[2637];
                        n_Body_y[2638] = c_Body_y[2637];
                    end else begin
                        n_Body_x[2638] = c_Body_x[c_Size-1];
                        n_Body_y[2638] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2639) begin
                        n_Body_x[2639] = c_Body_x[2638];
                        n_Body_y[2639] = c_Body_y[2638];
                    end else begin
                        n_Body_x[2639] = c_Body_x[c_Size-1];
                        n_Body_y[2639] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2640) begin
                        n_Body_x[2640] = c_Body_x[2639];
                        n_Body_y[2640] = c_Body_y[2639];
                    end else begin
                        n_Body_x[2640] = c_Body_x[c_Size-1];
                        n_Body_y[2640] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2641) begin
                        n_Body_x[2641] = c_Body_x[2640];
                        n_Body_y[2641] = c_Body_y[2640];
                    end else begin
                        n_Body_x[2641] = c_Body_x[c_Size-1];
                        n_Body_y[2641] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2642) begin
                        n_Body_x[2642] = c_Body_x[2641];
                        n_Body_y[2642] = c_Body_y[2641];
                    end else begin
                        n_Body_x[2642] = c_Body_x[c_Size-1];
                        n_Body_y[2642] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2643) begin
                        n_Body_x[2643] = c_Body_x[2642];
                        n_Body_y[2643] = c_Body_y[2642];
                    end else begin
                        n_Body_x[2643] = c_Body_x[c_Size-1];
                        n_Body_y[2643] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2644) begin
                        n_Body_x[2644] = c_Body_x[2643];
                        n_Body_y[2644] = c_Body_y[2643];
                    end else begin
                        n_Body_x[2644] = c_Body_x[c_Size-1];
                        n_Body_y[2644] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2645) begin
                        n_Body_x[2645] = c_Body_x[2644];
                        n_Body_y[2645] = c_Body_y[2644];
                    end else begin
                        n_Body_x[2645] = c_Body_x[c_Size-1];
                        n_Body_y[2645] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2646) begin
                        n_Body_x[2646] = c_Body_x[2645];
                        n_Body_y[2646] = c_Body_y[2645];
                    end else begin
                        n_Body_x[2646] = c_Body_x[c_Size-1];
                        n_Body_y[2646] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2647) begin
                        n_Body_x[2647] = c_Body_x[2646];
                        n_Body_y[2647] = c_Body_y[2646];
                    end else begin
                        n_Body_x[2647] = c_Body_x[c_Size-1];
                        n_Body_y[2647] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2648) begin
                        n_Body_x[2648] = c_Body_x[2647];
                        n_Body_y[2648] = c_Body_y[2647];
                    end else begin
                        n_Body_x[2648] = c_Body_x[c_Size-1];
                        n_Body_y[2648] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2649) begin
                        n_Body_x[2649] = c_Body_x[2648];
                        n_Body_y[2649] = c_Body_y[2648];
                    end else begin
                        n_Body_x[2649] = c_Body_x[c_Size-1];
                        n_Body_y[2649] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2650) begin
                        n_Body_x[2650] = c_Body_x[2649];
                        n_Body_y[2650] = c_Body_y[2649];
                    end else begin
                        n_Body_x[2650] = c_Body_x[c_Size-1];
                        n_Body_y[2650] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2651) begin
                        n_Body_x[2651] = c_Body_x[2650];
                        n_Body_y[2651] = c_Body_y[2650];
                    end else begin
                        n_Body_x[2651] = c_Body_x[c_Size-1];
                        n_Body_y[2651] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2652) begin
                        n_Body_x[2652] = c_Body_x[2651];
                        n_Body_y[2652] = c_Body_y[2651];
                    end else begin
                        n_Body_x[2652] = c_Body_x[c_Size-1];
                        n_Body_y[2652] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2653) begin
                        n_Body_x[2653] = c_Body_x[2652];
                        n_Body_y[2653] = c_Body_y[2652];
                    end else begin
                        n_Body_x[2653] = c_Body_x[c_Size-1];
                        n_Body_y[2653] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2654) begin
                        n_Body_x[2654] = c_Body_x[2653];
                        n_Body_y[2654] = c_Body_y[2653];
                    end else begin
                        n_Body_x[2654] = c_Body_x[c_Size-1];
                        n_Body_y[2654] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2655) begin
                        n_Body_x[2655] = c_Body_x[2654];
                        n_Body_y[2655] = c_Body_y[2654];
                    end else begin
                        n_Body_x[2655] = c_Body_x[c_Size-1];
                        n_Body_y[2655] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2656) begin
                        n_Body_x[2656] = c_Body_x[2655];
                        n_Body_y[2656] = c_Body_y[2655];
                    end else begin
                        n_Body_x[2656] = c_Body_x[c_Size-1];
                        n_Body_y[2656] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2657) begin
                        n_Body_x[2657] = c_Body_x[2656];
                        n_Body_y[2657] = c_Body_y[2656];
                    end else begin
                        n_Body_x[2657] = c_Body_x[c_Size-1];
                        n_Body_y[2657] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2658) begin
                        n_Body_x[2658] = c_Body_x[2657];
                        n_Body_y[2658] = c_Body_y[2657];
                    end else begin
                        n_Body_x[2658] = c_Body_x[c_Size-1];
                        n_Body_y[2658] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2659) begin
                        n_Body_x[2659] = c_Body_x[2658];
                        n_Body_y[2659] = c_Body_y[2658];
                    end else begin
                        n_Body_x[2659] = c_Body_x[c_Size-1];
                        n_Body_y[2659] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2660) begin
                        n_Body_x[2660] = c_Body_x[2659];
                        n_Body_y[2660] = c_Body_y[2659];
                    end else begin
                        n_Body_x[2660] = c_Body_x[c_Size-1];
                        n_Body_y[2660] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2661) begin
                        n_Body_x[2661] = c_Body_x[2660];
                        n_Body_y[2661] = c_Body_y[2660];
                    end else begin
                        n_Body_x[2661] = c_Body_x[c_Size-1];
                        n_Body_y[2661] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2662) begin
                        n_Body_x[2662] = c_Body_x[2661];
                        n_Body_y[2662] = c_Body_y[2661];
                    end else begin
                        n_Body_x[2662] = c_Body_x[c_Size-1];
                        n_Body_y[2662] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2663) begin
                        n_Body_x[2663] = c_Body_x[2662];
                        n_Body_y[2663] = c_Body_y[2662];
                    end else begin
                        n_Body_x[2663] = c_Body_x[c_Size-1];
                        n_Body_y[2663] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2664) begin
                        n_Body_x[2664] = c_Body_x[2663];
                        n_Body_y[2664] = c_Body_y[2663];
                    end else begin
                        n_Body_x[2664] = c_Body_x[c_Size-1];
                        n_Body_y[2664] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2665) begin
                        n_Body_x[2665] = c_Body_x[2664];
                        n_Body_y[2665] = c_Body_y[2664];
                    end else begin
                        n_Body_x[2665] = c_Body_x[c_Size-1];
                        n_Body_y[2665] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2666) begin
                        n_Body_x[2666] = c_Body_x[2665];
                        n_Body_y[2666] = c_Body_y[2665];
                    end else begin
                        n_Body_x[2666] = c_Body_x[c_Size-1];
                        n_Body_y[2666] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2667) begin
                        n_Body_x[2667] = c_Body_x[2666];
                        n_Body_y[2667] = c_Body_y[2666];
                    end else begin
                        n_Body_x[2667] = c_Body_x[c_Size-1];
                        n_Body_y[2667] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2668) begin
                        n_Body_x[2668] = c_Body_x[2667];
                        n_Body_y[2668] = c_Body_y[2667];
                    end else begin
                        n_Body_x[2668] = c_Body_x[c_Size-1];
                        n_Body_y[2668] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2669) begin
                        n_Body_x[2669] = c_Body_x[2668];
                        n_Body_y[2669] = c_Body_y[2668];
                    end else begin
                        n_Body_x[2669] = c_Body_x[c_Size-1];
                        n_Body_y[2669] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2670) begin
                        n_Body_x[2670] = c_Body_x[2669];
                        n_Body_y[2670] = c_Body_y[2669];
                    end else begin
                        n_Body_x[2670] = c_Body_x[c_Size-1];
                        n_Body_y[2670] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2671) begin
                        n_Body_x[2671] = c_Body_x[2670];
                        n_Body_y[2671] = c_Body_y[2670];
                    end else begin
                        n_Body_x[2671] = c_Body_x[c_Size-1];
                        n_Body_y[2671] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2672) begin
                        n_Body_x[2672] = c_Body_x[2671];
                        n_Body_y[2672] = c_Body_y[2671];
                    end else begin
                        n_Body_x[2672] = c_Body_x[c_Size-1];
                        n_Body_y[2672] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2673) begin
                        n_Body_x[2673] = c_Body_x[2672];
                        n_Body_y[2673] = c_Body_y[2672];
                    end else begin
                        n_Body_x[2673] = c_Body_x[c_Size-1];
                        n_Body_y[2673] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2674) begin
                        n_Body_x[2674] = c_Body_x[2673];
                        n_Body_y[2674] = c_Body_y[2673];
                    end else begin
                        n_Body_x[2674] = c_Body_x[c_Size-1];
                        n_Body_y[2674] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2675) begin
                        n_Body_x[2675] = c_Body_x[2674];
                        n_Body_y[2675] = c_Body_y[2674];
                    end else begin
                        n_Body_x[2675] = c_Body_x[c_Size-1];
                        n_Body_y[2675] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2676) begin
                        n_Body_x[2676] = c_Body_x[2675];
                        n_Body_y[2676] = c_Body_y[2675];
                    end else begin
                        n_Body_x[2676] = c_Body_x[c_Size-1];
                        n_Body_y[2676] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2677) begin
                        n_Body_x[2677] = c_Body_x[2676];
                        n_Body_y[2677] = c_Body_y[2676];
                    end else begin
                        n_Body_x[2677] = c_Body_x[c_Size-1];
                        n_Body_y[2677] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2678) begin
                        n_Body_x[2678] = c_Body_x[2677];
                        n_Body_y[2678] = c_Body_y[2677];
                    end else begin
                        n_Body_x[2678] = c_Body_x[c_Size-1];
                        n_Body_y[2678] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2679) begin
                        n_Body_x[2679] = c_Body_x[2678];
                        n_Body_y[2679] = c_Body_y[2678];
                    end else begin
                        n_Body_x[2679] = c_Body_x[c_Size-1];
                        n_Body_y[2679] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2680) begin
                        n_Body_x[2680] = c_Body_x[2679];
                        n_Body_y[2680] = c_Body_y[2679];
                    end else begin
                        n_Body_x[2680] = c_Body_x[c_Size-1];
                        n_Body_y[2680] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2681) begin
                        n_Body_x[2681] = c_Body_x[2680];
                        n_Body_y[2681] = c_Body_y[2680];
                    end else begin
                        n_Body_x[2681] = c_Body_x[c_Size-1];
                        n_Body_y[2681] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2682) begin
                        n_Body_x[2682] = c_Body_x[2681];
                        n_Body_y[2682] = c_Body_y[2681];
                    end else begin
                        n_Body_x[2682] = c_Body_x[c_Size-1];
                        n_Body_y[2682] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2683) begin
                        n_Body_x[2683] = c_Body_x[2682];
                        n_Body_y[2683] = c_Body_y[2682];
                    end else begin
                        n_Body_x[2683] = c_Body_x[c_Size-1];
                        n_Body_y[2683] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2684) begin
                        n_Body_x[2684] = c_Body_x[2683];
                        n_Body_y[2684] = c_Body_y[2683];
                    end else begin
                        n_Body_x[2684] = c_Body_x[c_Size-1];
                        n_Body_y[2684] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2685) begin
                        n_Body_x[2685] = c_Body_x[2684];
                        n_Body_y[2685] = c_Body_y[2684];
                    end else begin
                        n_Body_x[2685] = c_Body_x[c_Size-1];
                        n_Body_y[2685] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2686) begin
                        n_Body_x[2686] = c_Body_x[2685];
                        n_Body_y[2686] = c_Body_y[2685];
                    end else begin
                        n_Body_x[2686] = c_Body_x[c_Size-1];
                        n_Body_y[2686] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2687) begin
                        n_Body_x[2687] = c_Body_x[2686];
                        n_Body_y[2687] = c_Body_y[2686];
                    end else begin
                        n_Body_x[2687] = c_Body_x[c_Size-1];
                        n_Body_y[2687] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2688) begin
                        n_Body_x[2688] = c_Body_x[2687];
                        n_Body_y[2688] = c_Body_y[2687];
                    end else begin
                        n_Body_x[2688] = c_Body_x[c_Size-1];
                        n_Body_y[2688] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2689) begin
                        n_Body_x[2689] = c_Body_x[2688];
                        n_Body_y[2689] = c_Body_y[2688];
                    end else begin
                        n_Body_x[2689] = c_Body_x[c_Size-1];
                        n_Body_y[2689] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2690) begin
                        n_Body_x[2690] = c_Body_x[2689];
                        n_Body_y[2690] = c_Body_y[2689];
                    end else begin
                        n_Body_x[2690] = c_Body_x[c_Size-1];
                        n_Body_y[2690] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2691) begin
                        n_Body_x[2691] = c_Body_x[2690];
                        n_Body_y[2691] = c_Body_y[2690];
                    end else begin
                        n_Body_x[2691] = c_Body_x[c_Size-1];
                        n_Body_y[2691] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2692) begin
                        n_Body_x[2692] = c_Body_x[2691];
                        n_Body_y[2692] = c_Body_y[2691];
                    end else begin
                        n_Body_x[2692] = c_Body_x[c_Size-1];
                        n_Body_y[2692] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2693) begin
                        n_Body_x[2693] = c_Body_x[2692];
                        n_Body_y[2693] = c_Body_y[2692];
                    end else begin
                        n_Body_x[2693] = c_Body_x[c_Size-1];
                        n_Body_y[2693] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2694) begin
                        n_Body_x[2694] = c_Body_x[2693];
                        n_Body_y[2694] = c_Body_y[2693];
                    end else begin
                        n_Body_x[2694] = c_Body_x[c_Size-1];
                        n_Body_y[2694] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2695) begin
                        n_Body_x[2695] = c_Body_x[2694];
                        n_Body_y[2695] = c_Body_y[2694];
                    end else begin
                        n_Body_x[2695] = c_Body_x[c_Size-1];
                        n_Body_y[2695] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2696) begin
                        n_Body_x[2696] = c_Body_x[2695];
                        n_Body_y[2696] = c_Body_y[2695];
                    end else begin
                        n_Body_x[2696] = c_Body_x[c_Size-1];
                        n_Body_y[2696] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2697) begin
                        n_Body_x[2697] = c_Body_x[2696];
                        n_Body_y[2697] = c_Body_y[2696];
                    end else begin
                        n_Body_x[2697] = c_Body_x[c_Size-1];
                        n_Body_y[2697] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2698) begin
                        n_Body_x[2698] = c_Body_x[2697];
                        n_Body_y[2698] = c_Body_y[2697];
                    end else begin
                        n_Body_x[2698] = c_Body_x[c_Size-1];
                        n_Body_y[2698] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2699) begin
                        n_Body_x[2699] = c_Body_x[2698];
                        n_Body_y[2699] = c_Body_y[2698];
                    end else begin
                        n_Body_x[2699] = c_Body_x[c_Size-1];
                        n_Body_y[2699] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2700) begin
                        n_Body_x[2700] = c_Body_x[2699];
                        n_Body_y[2700] = c_Body_y[2699];
                    end else begin
                        n_Body_x[2700] = c_Body_x[c_Size-1];
                        n_Body_y[2700] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2701) begin
                        n_Body_x[2701] = c_Body_x[2700];
                        n_Body_y[2701] = c_Body_y[2700];
                    end else begin
                        n_Body_x[2701] = c_Body_x[c_Size-1];
                        n_Body_y[2701] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2702) begin
                        n_Body_x[2702] = c_Body_x[2701];
                        n_Body_y[2702] = c_Body_y[2701];
                    end else begin
                        n_Body_x[2702] = c_Body_x[c_Size-1];
                        n_Body_y[2702] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2703) begin
                        n_Body_x[2703] = c_Body_x[2702];
                        n_Body_y[2703] = c_Body_y[2702];
                    end else begin
                        n_Body_x[2703] = c_Body_x[c_Size-1];
                        n_Body_y[2703] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2704) begin
                        n_Body_x[2704] = c_Body_x[2703];
                        n_Body_y[2704] = c_Body_y[2703];
                    end else begin
                        n_Body_x[2704] = c_Body_x[c_Size-1];
                        n_Body_y[2704] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2705) begin
                        n_Body_x[2705] = c_Body_x[2704];
                        n_Body_y[2705] = c_Body_y[2704];
                    end else begin
                        n_Body_x[2705] = c_Body_x[c_Size-1];
                        n_Body_y[2705] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2706) begin
                        n_Body_x[2706] = c_Body_x[2705];
                        n_Body_y[2706] = c_Body_y[2705];
                    end else begin
                        n_Body_x[2706] = c_Body_x[c_Size-1];
                        n_Body_y[2706] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2707) begin
                        n_Body_x[2707] = c_Body_x[2706];
                        n_Body_y[2707] = c_Body_y[2706];
                    end else begin
                        n_Body_x[2707] = c_Body_x[c_Size-1];
                        n_Body_y[2707] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2708) begin
                        n_Body_x[2708] = c_Body_x[2707];
                        n_Body_y[2708] = c_Body_y[2707];
                    end else begin
                        n_Body_x[2708] = c_Body_x[c_Size-1];
                        n_Body_y[2708] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2709) begin
                        n_Body_x[2709] = c_Body_x[2708];
                        n_Body_y[2709] = c_Body_y[2708];
                    end else begin
                        n_Body_x[2709] = c_Body_x[c_Size-1];
                        n_Body_y[2709] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2710) begin
                        n_Body_x[2710] = c_Body_x[2709];
                        n_Body_y[2710] = c_Body_y[2709];
                    end else begin
                        n_Body_x[2710] = c_Body_x[c_Size-1];
                        n_Body_y[2710] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2711) begin
                        n_Body_x[2711] = c_Body_x[2710];
                        n_Body_y[2711] = c_Body_y[2710];
                    end else begin
                        n_Body_x[2711] = c_Body_x[c_Size-1];
                        n_Body_y[2711] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2712) begin
                        n_Body_x[2712] = c_Body_x[2711];
                        n_Body_y[2712] = c_Body_y[2711];
                    end else begin
                        n_Body_x[2712] = c_Body_x[c_Size-1];
                        n_Body_y[2712] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2713) begin
                        n_Body_x[2713] = c_Body_x[2712];
                        n_Body_y[2713] = c_Body_y[2712];
                    end else begin
                        n_Body_x[2713] = c_Body_x[c_Size-1];
                        n_Body_y[2713] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2714) begin
                        n_Body_x[2714] = c_Body_x[2713];
                        n_Body_y[2714] = c_Body_y[2713];
                    end else begin
                        n_Body_x[2714] = c_Body_x[c_Size-1];
                        n_Body_y[2714] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2715) begin
                        n_Body_x[2715] = c_Body_x[2714];
                        n_Body_y[2715] = c_Body_y[2714];
                    end else begin
                        n_Body_x[2715] = c_Body_x[c_Size-1];
                        n_Body_y[2715] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2716) begin
                        n_Body_x[2716] = c_Body_x[2715];
                        n_Body_y[2716] = c_Body_y[2715];
                    end else begin
                        n_Body_x[2716] = c_Body_x[c_Size-1];
                        n_Body_y[2716] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2717) begin
                        n_Body_x[2717] = c_Body_x[2716];
                        n_Body_y[2717] = c_Body_y[2716];
                    end else begin
                        n_Body_x[2717] = c_Body_x[c_Size-1];
                        n_Body_y[2717] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2718) begin
                        n_Body_x[2718] = c_Body_x[2717];
                        n_Body_y[2718] = c_Body_y[2717];
                    end else begin
                        n_Body_x[2718] = c_Body_x[c_Size-1];
                        n_Body_y[2718] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2719) begin
                        n_Body_x[2719] = c_Body_x[2718];
                        n_Body_y[2719] = c_Body_y[2718];
                    end else begin
                        n_Body_x[2719] = c_Body_x[c_Size-1];
                        n_Body_y[2719] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2720) begin
                        n_Body_x[2720] = c_Body_x[2719];
                        n_Body_y[2720] = c_Body_y[2719];
                    end else begin
                        n_Body_x[2720] = c_Body_x[c_Size-1];
                        n_Body_y[2720] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2721) begin
                        n_Body_x[2721] = c_Body_x[2720];
                        n_Body_y[2721] = c_Body_y[2720];
                    end else begin
                        n_Body_x[2721] = c_Body_x[c_Size-1];
                        n_Body_y[2721] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2722) begin
                        n_Body_x[2722] = c_Body_x[2721];
                        n_Body_y[2722] = c_Body_y[2721];
                    end else begin
                        n_Body_x[2722] = c_Body_x[c_Size-1];
                        n_Body_y[2722] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2723) begin
                        n_Body_x[2723] = c_Body_x[2722];
                        n_Body_y[2723] = c_Body_y[2722];
                    end else begin
                        n_Body_x[2723] = c_Body_x[c_Size-1];
                        n_Body_y[2723] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2724) begin
                        n_Body_x[2724] = c_Body_x[2723];
                        n_Body_y[2724] = c_Body_y[2723];
                    end else begin
                        n_Body_x[2724] = c_Body_x[c_Size-1];
                        n_Body_y[2724] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2725) begin
                        n_Body_x[2725] = c_Body_x[2724];
                        n_Body_y[2725] = c_Body_y[2724];
                    end else begin
                        n_Body_x[2725] = c_Body_x[c_Size-1];
                        n_Body_y[2725] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2726) begin
                        n_Body_x[2726] = c_Body_x[2725];
                        n_Body_y[2726] = c_Body_y[2725];
                    end else begin
                        n_Body_x[2726] = c_Body_x[c_Size-1];
                        n_Body_y[2726] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2727) begin
                        n_Body_x[2727] = c_Body_x[2726];
                        n_Body_y[2727] = c_Body_y[2726];
                    end else begin
                        n_Body_x[2727] = c_Body_x[c_Size-1];
                        n_Body_y[2727] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2728) begin
                        n_Body_x[2728] = c_Body_x[2727];
                        n_Body_y[2728] = c_Body_y[2727];
                    end else begin
                        n_Body_x[2728] = c_Body_x[c_Size-1];
                        n_Body_y[2728] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2729) begin
                        n_Body_x[2729] = c_Body_x[2728];
                        n_Body_y[2729] = c_Body_y[2728];
                    end else begin
                        n_Body_x[2729] = c_Body_x[c_Size-1];
                        n_Body_y[2729] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2730) begin
                        n_Body_x[2730] = c_Body_x[2729];
                        n_Body_y[2730] = c_Body_y[2729];
                    end else begin
                        n_Body_x[2730] = c_Body_x[c_Size-1];
                        n_Body_y[2730] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2731) begin
                        n_Body_x[2731] = c_Body_x[2730];
                        n_Body_y[2731] = c_Body_y[2730];
                    end else begin
                        n_Body_x[2731] = c_Body_x[c_Size-1];
                        n_Body_y[2731] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2732) begin
                        n_Body_x[2732] = c_Body_x[2731];
                        n_Body_y[2732] = c_Body_y[2731];
                    end else begin
                        n_Body_x[2732] = c_Body_x[c_Size-1];
                        n_Body_y[2732] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2733) begin
                        n_Body_x[2733] = c_Body_x[2732];
                        n_Body_y[2733] = c_Body_y[2732];
                    end else begin
                        n_Body_x[2733] = c_Body_x[c_Size-1];
                        n_Body_y[2733] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2734) begin
                        n_Body_x[2734] = c_Body_x[2733];
                        n_Body_y[2734] = c_Body_y[2733];
                    end else begin
                        n_Body_x[2734] = c_Body_x[c_Size-1];
                        n_Body_y[2734] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2735) begin
                        n_Body_x[2735] = c_Body_x[2734];
                        n_Body_y[2735] = c_Body_y[2734];
                    end else begin
                        n_Body_x[2735] = c_Body_x[c_Size-1];
                        n_Body_y[2735] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2736) begin
                        n_Body_x[2736] = c_Body_x[2735];
                        n_Body_y[2736] = c_Body_y[2735];
                    end else begin
                        n_Body_x[2736] = c_Body_x[c_Size-1];
                        n_Body_y[2736] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2737) begin
                        n_Body_x[2737] = c_Body_x[2736];
                        n_Body_y[2737] = c_Body_y[2736];
                    end else begin
                        n_Body_x[2737] = c_Body_x[c_Size-1];
                        n_Body_y[2737] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2738) begin
                        n_Body_x[2738] = c_Body_x[2737];
                        n_Body_y[2738] = c_Body_y[2737];
                    end else begin
                        n_Body_x[2738] = c_Body_x[c_Size-1];
                        n_Body_y[2738] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2739) begin
                        n_Body_x[2739] = c_Body_x[2738];
                        n_Body_y[2739] = c_Body_y[2738];
                    end else begin
                        n_Body_x[2739] = c_Body_x[c_Size-1];
                        n_Body_y[2739] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2740) begin
                        n_Body_x[2740] = c_Body_x[2739];
                        n_Body_y[2740] = c_Body_y[2739];
                    end else begin
                        n_Body_x[2740] = c_Body_x[c_Size-1];
                        n_Body_y[2740] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2741) begin
                        n_Body_x[2741] = c_Body_x[2740];
                        n_Body_y[2741] = c_Body_y[2740];
                    end else begin
                        n_Body_x[2741] = c_Body_x[c_Size-1];
                        n_Body_y[2741] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2742) begin
                        n_Body_x[2742] = c_Body_x[2741];
                        n_Body_y[2742] = c_Body_y[2741];
                    end else begin
                        n_Body_x[2742] = c_Body_x[c_Size-1];
                        n_Body_y[2742] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2743) begin
                        n_Body_x[2743] = c_Body_x[2742];
                        n_Body_y[2743] = c_Body_y[2742];
                    end else begin
                        n_Body_x[2743] = c_Body_x[c_Size-1];
                        n_Body_y[2743] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2744) begin
                        n_Body_x[2744] = c_Body_x[2743];
                        n_Body_y[2744] = c_Body_y[2743];
                    end else begin
                        n_Body_x[2744] = c_Body_x[c_Size-1];
                        n_Body_y[2744] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2745) begin
                        n_Body_x[2745] = c_Body_x[2744];
                        n_Body_y[2745] = c_Body_y[2744];
                    end else begin
                        n_Body_x[2745] = c_Body_x[c_Size-1];
                        n_Body_y[2745] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2746) begin
                        n_Body_x[2746] = c_Body_x[2745];
                        n_Body_y[2746] = c_Body_y[2745];
                    end else begin
                        n_Body_x[2746] = c_Body_x[c_Size-1];
                        n_Body_y[2746] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2747) begin
                        n_Body_x[2747] = c_Body_x[2746];
                        n_Body_y[2747] = c_Body_y[2746];
                    end else begin
                        n_Body_x[2747] = c_Body_x[c_Size-1];
                        n_Body_y[2747] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2748) begin
                        n_Body_x[2748] = c_Body_x[2747];
                        n_Body_y[2748] = c_Body_y[2747];
                    end else begin
                        n_Body_x[2748] = c_Body_x[c_Size-1];
                        n_Body_y[2748] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2749) begin
                        n_Body_x[2749] = c_Body_x[2748];
                        n_Body_y[2749] = c_Body_y[2748];
                    end else begin
                        n_Body_x[2749] = c_Body_x[c_Size-1];
                        n_Body_y[2749] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2750) begin
                        n_Body_x[2750] = c_Body_x[2749];
                        n_Body_y[2750] = c_Body_y[2749];
                    end else begin
                        n_Body_x[2750] = c_Body_x[c_Size-1];
                        n_Body_y[2750] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2751) begin
                        n_Body_x[2751] = c_Body_x[2750];
                        n_Body_y[2751] = c_Body_y[2750];
                    end else begin
                        n_Body_x[2751] = c_Body_x[c_Size-1];
                        n_Body_y[2751] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2752) begin
                        n_Body_x[2752] = c_Body_x[2751];
                        n_Body_y[2752] = c_Body_y[2751];
                    end else begin
                        n_Body_x[2752] = c_Body_x[c_Size-1];
                        n_Body_y[2752] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2753) begin
                        n_Body_x[2753] = c_Body_x[2752];
                        n_Body_y[2753] = c_Body_y[2752];
                    end else begin
                        n_Body_x[2753] = c_Body_x[c_Size-1];
                        n_Body_y[2753] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2754) begin
                        n_Body_x[2754] = c_Body_x[2753];
                        n_Body_y[2754] = c_Body_y[2753];
                    end else begin
                        n_Body_x[2754] = c_Body_x[c_Size-1];
                        n_Body_y[2754] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2755) begin
                        n_Body_x[2755] = c_Body_x[2754];
                        n_Body_y[2755] = c_Body_y[2754];
                    end else begin
                        n_Body_x[2755] = c_Body_x[c_Size-1];
                        n_Body_y[2755] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2756) begin
                        n_Body_x[2756] = c_Body_x[2755];
                        n_Body_y[2756] = c_Body_y[2755];
                    end else begin
                        n_Body_x[2756] = c_Body_x[c_Size-1];
                        n_Body_y[2756] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2757) begin
                        n_Body_x[2757] = c_Body_x[2756];
                        n_Body_y[2757] = c_Body_y[2756];
                    end else begin
                        n_Body_x[2757] = c_Body_x[c_Size-1];
                        n_Body_y[2757] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2758) begin
                        n_Body_x[2758] = c_Body_x[2757];
                        n_Body_y[2758] = c_Body_y[2757];
                    end else begin
                        n_Body_x[2758] = c_Body_x[c_Size-1];
                        n_Body_y[2758] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2759) begin
                        n_Body_x[2759] = c_Body_x[2758];
                        n_Body_y[2759] = c_Body_y[2758];
                    end else begin
                        n_Body_x[2759] = c_Body_x[c_Size-1];
                        n_Body_y[2759] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2760) begin
                        n_Body_x[2760] = c_Body_x[2759];
                        n_Body_y[2760] = c_Body_y[2759];
                    end else begin
                        n_Body_x[2760] = c_Body_x[c_Size-1];
                        n_Body_y[2760] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2761) begin
                        n_Body_x[2761] = c_Body_x[2760];
                        n_Body_y[2761] = c_Body_y[2760];
                    end else begin
                        n_Body_x[2761] = c_Body_x[c_Size-1];
                        n_Body_y[2761] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2762) begin
                        n_Body_x[2762] = c_Body_x[2761];
                        n_Body_y[2762] = c_Body_y[2761];
                    end else begin
                        n_Body_x[2762] = c_Body_x[c_Size-1];
                        n_Body_y[2762] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2763) begin
                        n_Body_x[2763] = c_Body_x[2762];
                        n_Body_y[2763] = c_Body_y[2762];
                    end else begin
                        n_Body_x[2763] = c_Body_x[c_Size-1];
                        n_Body_y[2763] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2764) begin
                        n_Body_x[2764] = c_Body_x[2763];
                        n_Body_y[2764] = c_Body_y[2763];
                    end else begin
                        n_Body_x[2764] = c_Body_x[c_Size-1];
                        n_Body_y[2764] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2765) begin
                        n_Body_x[2765] = c_Body_x[2764];
                        n_Body_y[2765] = c_Body_y[2764];
                    end else begin
                        n_Body_x[2765] = c_Body_x[c_Size-1];
                        n_Body_y[2765] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2766) begin
                        n_Body_x[2766] = c_Body_x[2765];
                        n_Body_y[2766] = c_Body_y[2765];
                    end else begin
                        n_Body_x[2766] = c_Body_x[c_Size-1];
                        n_Body_y[2766] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2767) begin
                        n_Body_x[2767] = c_Body_x[2766];
                        n_Body_y[2767] = c_Body_y[2766];
                    end else begin
                        n_Body_x[2767] = c_Body_x[c_Size-1];
                        n_Body_y[2767] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2768) begin
                        n_Body_x[2768] = c_Body_x[2767];
                        n_Body_y[2768] = c_Body_y[2767];
                    end else begin
                        n_Body_x[2768] = c_Body_x[c_Size-1];
                        n_Body_y[2768] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2769) begin
                        n_Body_x[2769] = c_Body_x[2768];
                        n_Body_y[2769] = c_Body_y[2768];
                    end else begin
                        n_Body_x[2769] = c_Body_x[c_Size-1];
                        n_Body_y[2769] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2770) begin
                        n_Body_x[2770] = c_Body_x[2769];
                        n_Body_y[2770] = c_Body_y[2769];
                    end else begin
                        n_Body_x[2770] = c_Body_x[c_Size-1];
                        n_Body_y[2770] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2771) begin
                        n_Body_x[2771] = c_Body_x[2770];
                        n_Body_y[2771] = c_Body_y[2770];
                    end else begin
                        n_Body_x[2771] = c_Body_x[c_Size-1];
                        n_Body_y[2771] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2772) begin
                        n_Body_x[2772] = c_Body_x[2771];
                        n_Body_y[2772] = c_Body_y[2771];
                    end else begin
                        n_Body_x[2772] = c_Body_x[c_Size-1];
                        n_Body_y[2772] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2773) begin
                        n_Body_x[2773] = c_Body_x[2772];
                        n_Body_y[2773] = c_Body_y[2772];
                    end else begin
                        n_Body_x[2773] = c_Body_x[c_Size-1];
                        n_Body_y[2773] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2774) begin
                        n_Body_x[2774] = c_Body_x[2773];
                        n_Body_y[2774] = c_Body_y[2773];
                    end else begin
                        n_Body_x[2774] = c_Body_x[c_Size-1];
                        n_Body_y[2774] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2775) begin
                        n_Body_x[2775] = c_Body_x[2774];
                        n_Body_y[2775] = c_Body_y[2774];
                    end else begin
                        n_Body_x[2775] = c_Body_x[c_Size-1];
                        n_Body_y[2775] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2776) begin
                        n_Body_x[2776] = c_Body_x[2775];
                        n_Body_y[2776] = c_Body_y[2775];
                    end else begin
                        n_Body_x[2776] = c_Body_x[c_Size-1];
                        n_Body_y[2776] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2777) begin
                        n_Body_x[2777] = c_Body_x[2776];
                        n_Body_y[2777] = c_Body_y[2776];
                    end else begin
                        n_Body_x[2777] = c_Body_x[c_Size-1];
                        n_Body_y[2777] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2778) begin
                        n_Body_x[2778] = c_Body_x[2777];
                        n_Body_y[2778] = c_Body_y[2777];
                    end else begin
                        n_Body_x[2778] = c_Body_x[c_Size-1];
                        n_Body_y[2778] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2779) begin
                        n_Body_x[2779] = c_Body_x[2778];
                        n_Body_y[2779] = c_Body_y[2778];
                    end else begin
                        n_Body_x[2779] = c_Body_x[c_Size-1];
                        n_Body_y[2779] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2780) begin
                        n_Body_x[2780] = c_Body_x[2779];
                        n_Body_y[2780] = c_Body_y[2779];
                    end else begin
                        n_Body_x[2780] = c_Body_x[c_Size-1];
                        n_Body_y[2780] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2781) begin
                        n_Body_x[2781] = c_Body_x[2780];
                        n_Body_y[2781] = c_Body_y[2780];
                    end else begin
                        n_Body_x[2781] = c_Body_x[c_Size-1];
                        n_Body_y[2781] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2782) begin
                        n_Body_x[2782] = c_Body_x[2781];
                        n_Body_y[2782] = c_Body_y[2781];
                    end else begin
                        n_Body_x[2782] = c_Body_x[c_Size-1];
                        n_Body_y[2782] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2783) begin
                        n_Body_x[2783] = c_Body_x[2782];
                        n_Body_y[2783] = c_Body_y[2782];
                    end else begin
                        n_Body_x[2783] = c_Body_x[c_Size-1];
                        n_Body_y[2783] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2784) begin
                        n_Body_x[2784] = c_Body_x[2783];
                        n_Body_y[2784] = c_Body_y[2783];
                    end else begin
                        n_Body_x[2784] = c_Body_x[c_Size-1];
                        n_Body_y[2784] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2785) begin
                        n_Body_x[2785] = c_Body_x[2784];
                        n_Body_y[2785] = c_Body_y[2784];
                    end else begin
                        n_Body_x[2785] = c_Body_x[c_Size-1];
                        n_Body_y[2785] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2786) begin
                        n_Body_x[2786] = c_Body_x[2785];
                        n_Body_y[2786] = c_Body_y[2785];
                    end else begin
                        n_Body_x[2786] = c_Body_x[c_Size-1];
                        n_Body_y[2786] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2787) begin
                        n_Body_x[2787] = c_Body_x[2786];
                        n_Body_y[2787] = c_Body_y[2786];
                    end else begin
                        n_Body_x[2787] = c_Body_x[c_Size-1];
                        n_Body_y[2787] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2788) begin
                        n_Body_x[2788] = c_Body_x[2787];
                        n_Body_y[2788] = c_Body_y[2787];
                    end else begin
                        n_Body_x[2788] = c_Body_x[c_Size-1];
                        n_Body_y[2788] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2789) begin
                        n_Body_x[2789] = c_Body_x[2788];
                        n_Body_y[2789] = c_Body_y[2788];
                    end else begin
                        n_Body_x[2789] = c_Body_x[c_Size-1];
                        n_Body_y[2789] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2790) begin
                        n_Body_x[2790] = c_Body_x[2789];
                        n_Body_y[2790] = c_Body_y[2789];
                    end else begin
                        n_Body_x[2790] = c_Body_x[c_Size-1];
                        n_Body_y[2790] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2791) begin
                        n_Body_x[2791] = c_Body_x[2790];
                        n_Body_y[2791] = c_Body_y[2790];
                    end else begin
                        n_Body_x[2791] = c_Body_x[c_Size-1];
                        n_Body_y[2791] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2792) begin
                        n_Body_x[2792] = c_Body_x[2791];
                        n_Body_y[2792] = c_Body_y[2791];
                    end else begin
                        n_Body_x[2792] = c_Body_x[c_Size-1];
                        n_Body_y[2792] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2793) begin
                        n_Body_x[2793] = c_Body_x[2792];
                        n_Body_y[2793] = c_Body_y[2792];
                    end else begin
                        n_Body_x[2793] = c_Body_x[c_Size-1];
                        n_Body_y[2793] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2794) begin
                        n_Body_x[2794] = c_Body_x[2793];
                        n_Body_y[2794] = c_Body_y[2793];
                    end else begin
                        n_Body_x[2794] = c_Body_x[c_Size-1];
                        n_Body_y[2794] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2795) begin
                        n_Body_x[2795] = c_Body_x[2794];
                        n_Body_y[2795] = c_Body_y[2794];
                    end else begin
                        n_Body_x[2795] = c_Body_x[c_Size-1];
                        n_Body_y[2795] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2796) begin
                        n_Body_x[2796] = c_Body_x[2795];
                        n_Body_y[2796] = c_Body_y[2795];
                    end else begin
                        n_Body_x[2796] = c_Body_x[c_Size-1];
                        n_Body_y[2796] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2797) begin
                        n_Body_x[2797] = c_Body_x[2796];
                        n_Body_y[2797] = c_Body_y[2796];
                    end else begin
                        n_Body_x[2797] = c_Body_x[c_Size-1];
                        n_Body_y[2797] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2798) begin
                        n_Body_x[2798] = c_Body_x[2797];
                        n_Body_y[2798] = c_Body_y[2797];
                    end else begin
                        n_Body_x[2798] = c_Body_x[c_Size-1];
                        n_Body_y[2798] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2799) begin
                        n_Body_x[2799] = c_Body_x[2798];
                        n_Body_y[2799] = c_Body_y[2798];
                    end else begin
                        n_Body_x[2799] = c_Body_x[c_Size-1];
                        n_Body_y[2799] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2800) begin
                        n_Body_x[2800] = c_Body_x[2799];
                        n_Body_y[2800] = c_Body_y[2799];
                    end else begin
                        n_Body_x[2800] = c_Body_x[c_Size-1];
                        n_Body_y[2800] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2801) begin
                        n_Body_x[2801] = c_Body_x[2800];
                        n_Body_y[2801] = c_Body_y[2800];
                    end else begin
                        n_Body_x[2801] = c_Body_x[c_Size-1];
                        n_Body_y[2801] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2802) begin
                        n_Body_x[2802] = c_Body_x[2801];
                        n_Body_y[2802] = c_Body_y[2801];
                    end else begin
                        n_Body_x[2802] = c_Body_x[c_Size-1];
                        n_Body_y[2802] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2803) begin
                        n_Body_x[2803] = c_Body_x[2802];
                        n_Body_y[2803] = c_Body_y[2802];
                    end else begin
                        n_Body_x[2803] = c_Body_x[c_Size-1];
                        n_Body_y[2803] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2804) begin
                        n_Body_x[2804] = c_Body_x[2803];
                        n_Body_y[2804] = c_Body_y[2803];
                    end else begin
                        n_Body_x[2804] = c_Body_x[c_Size-1];
                        n_Body_y[2804] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2805) begin
                        n_Body_x[2805] = c_Body_x[2804];
                        n_Body_y[2805] = c_Body_y[2804];
                    end else begin
                        n_Body_x[2805] = c_Body_x[c_Size-1];
                        n_Body_y[2805] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2806) begin
                        n_Body_x[2806] = c_Body_x[2805];
                        n_Body_y[2806] = c_Body_y[2805];
                    end else begin
                        n_Body_x[2806] = c_Body_x[c_Size-1];
                        n_Body_y[2806] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2807) begin
                        n_Body_x[2807] = c_Body_x[2806];
                        n_Body_y[2807] = c_Body_y[2806];
                    end else begin
                        n_Body_x[2807] = c_Body_x[c_Size-1];
                        n_Body_y[2807] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2808) begin
                        n_Body_x[2808] = c_Body_x[2807];
                        n_Body_y[2808] = c_Body_y[2807];
                    end else begin
                        n_Body_x[2808] = c_Body_x[c_Size-1];
                        n_Body_y[2808] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2809) begin
                        n_Body_x[2809] = c_Body_x[2808];
                        n_Body_y[2809] = c_Body_y[2808];
                    end else begin
                        n_Body_x[2809] = c_Body_x[c_Size-1];
                        n_Body_y[2809] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2810) begin
                        n_Body_x[2810] = c_Body_x[2809];
                        n_Body_y[2810] = c_Body_y[2809];
                    end else begin
                        n_Body_x[2810] = c_Body_x[c_Size-1];
                        n_Body_y[2810] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2811) begin
                        n_Body_x[2811] = c_Body_x[2810];
                        n_Body_y[2811] = c_Body_y[2810];
                    end else begin
                        n_Body_x[2811] = c_Body_x[c_Size-1];
                        n_Body_y[2811] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2812) begin
                        n_Body_x[2812] = c_Body_x[2811];
                        n_Body_y[2812] = c_Body_y[2811];
                    end else begin
                        n_Body_x[2812] = c_Body_x[c_Size-1];
                        n_Body_y[2812] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2813) begin
                        n_Body_x[2813] = c_Body_x[2812];
                        n_Body_y[2813] = c_Body_y[2812];
                    end else begin
                        n_Body_x[2813] = c_Body_x[c_Size-1];
                        n_Body_y[2813] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2814) begin
                        n_Body_x[2814] = c_Body_x[2813];
                        n_Body_y[2814] = c_Body_y[2813];
                    end else begin
                        n_Body_x[2814] = c_Body_x[c_Size-1];
                        n_Body_y[2814] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2815) begin
                        n_Body_x[2815] = c_Body_x[2814];
                        n_Body_y[2815] = c_Body_y[2814];
                    end else begin
                        n_Body_x[2815] = c_Body_x[c_Size-1];
                        n_Body_y[2815] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2816) begin
                        n_Body_x[2816] = c_Body_x[2815];
                        n_Body_y[2816] = c_Body_y[2815];
                    end else begin
                        n_Body_x[2816] = c_Body_x[c_Size-1];
                        n_Body_y[2816] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2817) begin
                        n_Body_x[2817] = c_Body_x[2816];
                        n_Body_y[2817] = c_Body_y[2816];
                    end else begin
                        n_Body_x[2817] = c_Body_x[c_Size-1];
                        n_Body_y[2817] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2818) begin
                        n_Body_x[2818] = c_Body_x[2817];
                        n_Body_y[2818] = c_Body_y[2817];
                    end else begin
                        n_Body_x[2818] = c_Body_x[c_Size-1];
                        n_Body_y[2818] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2819) begin
                        n_Body_x[2819] = c_Body_x[2818];
                        n_Body_y[2819] = c_Body_y[2818];
                    end else begin
                        n_Body_x[2819] = c_Body_x[c_Size-1];
                        n_Body_y[2819] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2820) begin
                        n_Body_x[2820] = c_Body_x[2819];
                        n_Body_y[2820] = c_Body_y[2819];
                    end else begin
                        n_Body_x[2820] = c_Body_x[c_Size-1];
                        n_Body_y[2820] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2821) begin
                        n_Body_x[2821] = c_Body_x[2820];
                        n_Body_y[2821] = c_Body_y[2820];
                    end else begin
                        n_Body_x[2821] = c_Body_x[c_Size-1];
                        n_Body_y[2821] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2822) begin
                        n_Body_x[2822] = c_Body_x[2821];
                        n_Body_y[2822] = c_Body_y[2821];
                    end else begin
                        n_Body_x[2822] = c_Body_x[c_Size-1];
                        n_Body_y[2822] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2823) begin
                        n_Body_x[2823] = c_Body_x[2822];
                        n_Body_y[2823] = c_Body_y[2822];
                    end else begin
                        n_Body_x[2823] = c_Body_x[c_Size-1];
                        n_Body_y[2823] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2824) begin
                        n_Body_x[2824] = c_Body_x[2823];
                        n_Body_y[2824] = c_Body_y[2823];
                    end else begin
                        n_Body_x[2824] = c_Body_x[c_Size-1];
                        n_Body_y[2824] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2825) begin
                        n_Body_x[2825] = c_Body_x[2824];
                        n_Body_y[2825] = c_Body_y[2824];
                    end else begin
                        n_Body_x[2825] = c_Body_x[c_Size-1];
                        n_Body_y[2825] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2826) begin
                        n_Body_x[2826] = c_Body_x[2825];
                        n_Body_y[2826] = c_Body_y[2825];
                    end else begin
                        n_Body_x[2826] = c_Body_x[c_Size-1];
                        n_Body_y[2826] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2827) begin
                        n_Body_x[2827] = c_Body_x[2826];
                        n_Body_y[2827] = c_Body_y[2826];
                    end else begin
                        n_Body_x[2827] = c_Body_x[c_Size-1];
                        n_Body_y[2827] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2828) begin
                        n_Body_x[2828] = c_Body_x[2827];
                        n_Body_y[2828] = c_Body_y[2827];
                    end else begin
                        n_Body_x[2828] = c_Body_x[c_Size-1];
                        n_Body_y[2828] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2829) begin
                        n_Body_x[2829] = c_Body_x[2828];
                        n_Body_y[2829] = c_Body_y[2828];
                    end else begin
                        n_Body_x[2829] = c_Body_x[c_Size-1];
                        n_Body_y[2829] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2830) begin
                        n_Body_x[2830] = c_Body_x[2829];
                        n_Body_y[2830] = c_Body_y[2829];
                    end else begin
                        n_Body_x[2830] = c_Body_x[c_Size-1];
                        n_Body_y[2830] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2831) begin
                        n_Body_x[2831] = c_Body_x[2830];
                        n_Body_y[2831] = c_Body_y[2830];
                    end else begin
                        n_Body_x[2831] = c_Body_x[c_Size-1];
                        n_Body_y[2831] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2832) begin
                        n_Body_x[2832] = c_Body_x[2831];
                        n_Body_y[2832] = c_Body_y[2831];
                    end else begin
                        n_Body_x[2832] = c_Body_x[c_Size-1];
                        n_Body_y[2832] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2833) begin
                        n_Body_x[2833] = c_Body_x[2832];
                        n_Body_y[2833] = c_Body_y[2832];
                    end else begin
                        n_Body_x[2833] = c_Body_x[c_Size-1];
                        n_Body_y[2833] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2834) begin
                        n_Body_x[2834] = c_Body_x[2833];
                        n_Body_y[2834] = c_Body_y[2833];
                    end else begin
                        n_Body_x[2834] = c_Body_x[c_Size-1];
                        n_Body_y[2834] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2835) begin
                        n_Body_x[2835] = c_Body_x[2834];
                        n_Body_y[2835] = c_Body_y[2834];
                    end else begin
                        n_Body_x[2835] = c_Body_x[c_Size-1];
                        n_Body_y[2835] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2836) begin
                        n_Body_x[2836] = c_Body_x[2835];
                        n_Body_y[2836] = c_Body_y[2835];
                    end else begin
                        n_Body_x[2836] = c_Body_x[c_Size-1];
                        n_Body_y[2836] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2837) begin
                        n_Body_x[2837] = c_Body_x[2836];
                        n_Body_y[2837] = c_Body_y[2836];
                    end else begin
                        n_Body_x[2837] = c_Body_x[c_Size-1];
                        n_Body_y[2837] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2838) begin
                        n_Body_x[2838] = c_Body_x[2837];
                        n_Body_y[2838] = c_Body_y[2837];
                    end else begin
                        n_Body_x[2838] = c_Body_x[c_Size-1];
                        n_Body_y[2838] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2839) begin
                        n_Body_x[2839] = c_Body_x[2838];
                        n_Body_y[2839] = c_Body_y[2838];
                    end else begin
                        n_Body_x[2839] = c_Body_x[c_Size-1];
                        n_Body_y[2839] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2840) begin
                        n_Body_x[2840] = c_Body_x[2839];
                        n_Body_y[2840] = c_Body_y[2839];
                    end else begin
                        n_Body_x[2840] = c_Body_x[c_Size-1];
                        n_Body_y[2840] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2841) begin
                        n_Body_x[2841] = c_Body_x[2840];
                        n_Body_y[2841] = c_Body_y[2840];
                    end else begin
                        n_Body_x[2841] = c_Body_x[c_Size-1];
                        n_Body_y[2841] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2842) begin
                        n_Body_x[2842] = c_Body_x[2841];
                        n_Body_y[2842] = c_Body_y[2841];
                    end else begin
                        n_Body_x[2842] = c_Body_x[c_Size-1];
                        n_Body_y[2842] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2843) begin
                        n_Body_x[2843] = c_Body_x[2842];
                        n_Body_y[2843] = c_Body_y[2842];
                    end else begin
                        n_Body_x[2843] = c_Body_x[c_Size-1];
                        n_Body_y[2843] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2844) begin
                        n_Body_x[2844] = c_Body_x[2843];
                        n_Body_y[2844] = c_Body_y[2843];
                    end else begin
                        n_Body_x[2844] = c_Body_x[c_Size-1];
                        n_Body_y[2844] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2845) begin
                        n_Body_x[2845] = c_Body_x[2844];
                        n_Body_y[2845] = c_Body_y[2844];
                    end else begin
                        n_Body_x[2845] = c_Body_x[c_Size-1];
                        n_Body_y[2845] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2846) begin
                        n_Body_x[2846] = c_Body_x[2845];
                        n_Body_y[2846] = c_Body_y[2845];
                    end else begin
                        n_Body_x[2846] = c_Body_x[c_Size-1];
                        n_Body_y[2846] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2847) begin
                        n_Body_x[2847] = c_Body_x[2846];
                        n_Body_y[2847] = c_Body_y[2846];
                    end else begin
                        n_Body_x[2847] = c_Body_x[c_Size-1];
                        n_Body_y[2847] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2848) begin
                        n_Body_x[2848] = c_Body_x[2847];
                        n_Body_y[2848] = c_Body_y[2847];
                    end else begin
                        n_Body_x[2848] = c_Body_x[c_Size-1];
                        n_Body_y[2848] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2849) begin
                        n_Body_x[2849] = c_Body_x[2848];
                        n_Body_y[2849] = c_Body_y[2848];
                    end else begin
                        n_Body_x[2849] = c_Body_x[c_Size-1];
                        n_Body_y[2849] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2850) begin
                        n_Body_x[2850] = c_Body_x[2849];
                        n_Body_y[2850] = c_Body_y[2849];
                    end else begin
                        n_Body_x[2850] = c_Body_x[c_Size-1];
                        n_Body_y[2850] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2851) begin
                        n_Body_x[2851] = c_Body_x[2850];
                        n_Body_y[2851] = c_Body_y[2850];
                    end else begin
                        n_Body_x[2851] = c_Body_x[c_Size-1];
                        n_Body_y[2851] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2852) begin
                        n_Body_x[2852] = c_Body_x[2851];
                        n_Body_y[2852] = c_Body_y[2851];
                    end else begin
                        n_Body_x[2852] = c_Body_x[c_Size-1];
                        n_Body_y[2852] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2853) begin
                        n_Body_x[2853] = c_Body_x[2852];
                        n_Body_y[2853] = c_Body_y[2852];
                    end else begin
                        n_Body_x[2853] = c_Body_x[c_Size-1];
                        n_Body_y[2853] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2854) begin
                        n_Body_x[2854] = c_Body_x[2853];
                        n_Body_y[2854] = c_Body_y[2853];
                    end else begin
                        n_Body_x[2854] = c_Body_x[c_Size-1];
                        n_Body_y[2854] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2855) begin
                        n_Body_x[2855] = c_Body_x[2854];
                        n_Body_y[2855] = c_Body_y[2854];
                    end else begin
                        n_Body_x[2855] = c_Body_x[c_Size-1];
                        n_Body_y[2855] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2856) begin
                        n_Body_x[2856] = c_Body_x[2855];
                        n_Body_y[2856] = c_Body_y[2855];
                    end else begin
                        n_Body_x[2856] = c_Body_x[c_Size-1];
                        n_Body_y[2856] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2857) begin
                        n_Body_x[2857] = c_Body_x[2856];
                        n_Body_y[2857] = c_Body_y[2856];
                    end else begin
                        n_Body_x[2857] = c_Body_x[c_Size-1];
                        n_Body_y[2857] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2858) begin
                        n_Body_x[2858] = c_Body_x[2857];
                        n_Body_y[2858] = c_Body_y[2857];
                    end else begin
                        n_Body_x[2858] = c_Body_x[c_Size-1];
                        n_Body_y[2858] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2859) begin
                        n_Body_x[2859] = c_Body_x[2858];
                        n_Body_y[2859] = c_Body_y[2858];
                    end else begin
                        n_Body_x[2859] = c_Body_x[c_Size-1];
                        n_Body_y[2859] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2860) begin
                        n_Body_x[2860] = c_Body_x[2859];
                        n_Body_y[2860] = c_Body_y[2859];
                    end else begin
                        n_Body_x[2860] = c_Body_x[c_Size-1];
                        n_Body_y[2860] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2861) begin
                        n_Body_x[2861] = c_Body_x[2860];
                        n_Body_y[2861] = c_Body_y[2860];
                    end else begin
                        n_Body_x[2861] = c_Body_x[c_Size-1];
                        n_Body_y[2861] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2862) begin
                        n_Body_x[2862] = c_Body_x[2861];
                        n_Body_y[2862] = c_Body_y[2861];
                    end else begin
                        n_Body_x[2862] = c_Body_x[c_Size-1];
                        n_Body_y[2862] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2863) begin
                        n_Body_x[2863] = c_Body_x[2862];
                        n_Body_y[2863] = c_Body_y[2862];
                    end else begin
                        n_Body_x[2863] = c_Body_x[c_Size-1];
                        n_Body_y[2863] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2864) begin
                        n_Body_x[2864] = c_Body_x[2863];
                        n_Body_y[2864] = c_Body_y[2863];
                    end else begin
                        n_Body_x[2864] = c_Body_x[c_Size-1];
                        n_Body_y[2864] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2865) begin
                        n_Body_x[2865] = c_Body_x[2864];
                        n_Body_y[2865] = c_Body_y[2864];
                    end else begin
                        n_Body_x[2865] = c_Body_x[c_Size-1];
                        n_Body_y[2865] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2866) begin
                        n_Body_x[2866] = c_Body_x[2865];
                        n_Body_y[2866] = c_Body_y[2865];
                    end else begin
                        n_Body_x[2866] = c_Body_x[c_Size-1];
                        n_Body_y[2866] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2867) begin
                        n_Body_x[2867] = c_Body_x[2866];
                        n_Body_y[2867] = c_Body_y[2866];
                    end else begin
                        n_Body_x[2867] = c_Body_x[c_Size-1];
                        n_Body_y[2867] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2868) begin
                        n_Body_x[2868] = c_Body_x[2867];
                        n_Body_y[2868] = c_Body_y[2867];
                    end else begin
                        n_Body_x[2868] = c_Body_x[c_Size-1];
                        n_Body_y[2868] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2869) begin
                        n_Body_x[2869] = c_Body_x[2868];
                        n_Body_y[2869] = c_Body_y[2868];
                    end else begin
                        n_Body_x[2869] = c_Body_x[c_Size-1];
                        n_Body_y[2869] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2870) begin
                        n_Body_x[2870] = c_Body_x[2869];
                        n_Body_y[2870] = c_Body_y[2869];
                    end else begin
                        n_Body_x[2870] = c_Body_x[c_Size-1];
                        n_Body_y[2870] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2871) begin
                        n_Body_x[2871] = c_Body_x[2870];
                        n_Body_y[2871] = c_Body_y[2870];
                    end else begin
                        n_Body_x[2871] = c_Body_x[c_Size-1];
                        n_Body_y[2871] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2872) begin
                        n_Body_x[2872] = c_Body_x[2871];
                        n_Body_y[2872] = c_Body_y[2871];
                    end else begin
                        n_Body_x[2872] = c_Body_x[c_Size-1];
                        n_Body_y[2872] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2873) begin
                        n_Body_x[2873] = c_Body_x[2872];
                        n_Body_y[2873] = c_Body_y[2872];
                    end else begin
                        n_Body_x[2873] = c_Body_x[c_Size-1];
                        n_Body_y[2873] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2874) begin
                        n_Body_x[2874] = c_Body_x[2873];
                        n_Body_y[2874] = c_Body_y[2873];
                    end else begin
                        n_Body_x[2874] = c_Body_x[c_Size-1];
                        n_Body_y[2874] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2875) begin
                        n_Body_x[2875] = c_Body_x[2874];
                        n_Body_y[2875] = c_Body_y[2874];
                    end else begin
                        n_Body_x[2875] = c_Body_x[c_Size-1];
                        n_Body_y[2875] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2876) begin
                        n_Body_x[2876] = c_Body_x[2875];
                        n_Body_y[2876] = c_Body_y[2875];
                    end else begin
                        n_Body_x[2876] = c_Body_x[c_Size-1];
                        n_Body_y[2876] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2877) begin
                        n_Body_x[2877] = c_Body_x[2876];
                        n_Body_y[2877] = c_Body_y[2876];
                    end else begin
                        n_Body_x[2877] = c_Body_x[c_Size-1];
                        n_Body_y[2877] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2878) begin
                        n_Body_x[2878] = c_Body_x[2877];
                        n_Body_y[2878] = c_Body_y[2877];
                    end else begin
                        n_Body_x[2878] = c_Body_x[c_Size-1];
                        n_Body_y[2878] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2879) begin
                        n_Body_x[2879] = c_Body_x[2878];
                        n_Body_y[2879] = c_Body_y[2878];
                    end else begin
                        n_Body_x[2879] = c_Body_x[c_Size-1];
                        n_Body_y[2879] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2880) begin
                        n_Body_x[2880] = c_Body_x[2879];
                        n_Body_y[2880] = c_Body_y[2879];
                    end else begin
                        n_Body_x[2880] = c_Body_x[c_Size-1];
                        n_Body_y[2880] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2881) begin
                        n_Body_x[2881] = c_Body_x[2880];
                        n_Body_y[2881] = c_Body_y[2880];
                    end else begin
                        n_Body_x[2881] = c_Body_x[c_Size-1];
                        n_Body_y[2881] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2882) begin
                        n_Body_x[2882] = c_Body_x[2881];
                        n_Body_y[2882] = c_Body_y[2881];
                    end else begin
                        n_Body_x[2882] = c_Body_x[c_Size-1];
                        n_Body_y[2882] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2883) begin
                        n_Body_x[2883] = c_Body_x[2882];
                        n_Body_y[2883] = c_Body_y[2882];
                    end else begin
                        n_Body_x[2883] = c_Body_x[c_Size-1];
                        n_Body_y[2883] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2884) begin
                        n_Body_x[2884] = c_Body_x[2883];
                        n_Body_y[2884] = c_Body_y[2883];
                    end else begin
                        n_Body_x[2884] = c_Body_x[c_Size-1];
                        n_Body_y[2884] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2885) begin
                        n_Body_x[2885] = c_Body_x[2884];
                        n_Body_y[2885] = c_Body_y[2884];
                    end else begin
                        n_Body_x[2885] = c_Body_x[c_Size-1];
                        n_Body_y[2885] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2886) begin
                        n_Body_x[2886] = c_Body_x[2885];
                        n_Body_y[2886] = c_Body_y[2885];
                    end else begin
                        n_Body_x[2886] = c_Body_x[c_Size-1];
                        n_Body_y[2886] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2887) begin
                        n_Body_x[2887] = c_Body_x[2886];
                        n_Body_y[2887] = c_Body_y[2886];
                    end else begin
                        n_Body_x[2887] = c_Body_x[c_Size-1];
                        n_Body_y[2887] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2888) begin
                        n_Body_x[2888] = c_Body_x[2887];
                        n_Body_y[2888] = c_Body_y[2887];
                    end else begin
                        n_Body_x[2888] = c_Body_x[c_Size-1];
                        n_Body_y[2888] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2889) begin
                        n_Body_x[2889] = c_Body_x[2888];
                        n_Body_y[2889] = c_Body_y[2888];
                    end else begin
                        n_Body_x[2889] = c_Body_x[c_Size-1];
                        n_Body_y[2889] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2890) begin
                        n_Body_x[2890] = c_Body_x[2889];
                        n_Body_y[2890] = c_Body_y[2889];
                    end else begin
                        n_Body_x[2890] = c_Body_x[c_Size-1];
                        n_Body_y[2890] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2891) begin
                        n_Body_x[2891] = c_Body_x[2890];
                        n_Body_y[2891] = c_Body_y[2890];
                    end else begin
                        n_Body_x[2891] = c_Body_x[c_Size-1];
                        n_Body_y[2891] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2892) begin
                        n_Body_x[2892] = c_Body_x[2891];
                        n_Body_y[2892] = c_Body_y[2891];
                    end else begin
                        n_Body_x[2892] = c_Body_x[c_Size-1];
                        n_Body_y[2892] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2893) begin
                        n_Body_x[2893] = c_Body_x[2892];
                        n_Body_y[2893] = c_Body_y[2892];
                    end else begin
                        n_Body_x[2893] = c_Body_x[c_Size-1];
                        n_Body_y[2893] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2894) begin
                        n_Body_x[2894] = c_Body_x[2893];
                        n_Body_y[2894] = c_Body_y[2893];
                    end else begin
                        n_Body_x[2894] = c_Body_x[c_Size-1];
                        n_Body_y[2894] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2895) begin
                        n_Body_x[2895] = c_Body_x[2894];
                        n_Body_y[2895] = c_Body_y[2894];
                    end else begin
                        n_Body_x[2895] = c_Body_x[c_Size-1];
                        n_Body_y[2895] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2896) begin
                        n_Body_x[2896] = c_Body_x[2895];
                        n_Body_y[2896] = c_Body_y[2895];
                    end else begin
                        n_Body_x[2896] = c_Body_x[c_Size-1];
                        n_Body_y[2896] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2897) begin
                        n_Body_x[2897] = c_Body_x[2896];
                        n_Body_y[2897] = c_Body_y[2896];
                    end else begin
                        n_Body_x[2897] = c_Body_x[c_Size-1];
                        n_Body_y[2897] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2898) begin
                        n_Body_x[2898] = c_Body_x[2897];
                        n_Body_y[2898] = c_Body_y[2897];
                    end else begin
                        n_Body_x[2898] = c_Body_x[c_Size-1];
                        n_Body_y[2898] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2899) begin
                        n_Body_x[2899] = c_Body_x[2898];
                        n_Body_y[2899] = c_Body_y[2898];
                    end else begin
                        n_Body_x[2899] = c_Body_x[c_Size-1];
                        n_Body_y[2899] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2900) begin
                        n_Body_x[2900] = c_Body_x[2899];
                        n_Body_y[2900] = c_Body_y[2899];
                    end else begin
                        n_Body_x[2900] = c_Body_x[c_Size-1];
                        n_Body_y[2900] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2901) begin
                        n_Body_x[2901] = c_Body_x[2900];
                        n_Body_y[2901] = c_Body_y[2900];
                    end else begin
                        n_Body_x[2901] = c_Body_x[c_Size-1];
                        n_Body_y[2901] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2902) begin
                        n_Body_x[2902] = c_Body_x[2901];
                        n_Body_y[2902] = c_Body_y[2901];
                    end else begin
                        n_Body_x[2902] = c_Body_x[c_Size-1];
                        n_Body_y[2902] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2903) begin
                        n_Body_x[2903] = c_Body_x[2902];
                        n_Body_y[2903] = c_Body_y[2902];
                    end else begin
                        n_Body_x[2903] = c_Body_x[c_Size-1];
                        n_Body_y[2903] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2904) begin
                        n_Body_x[2904] = c_Body_x[2903];
                        n_Body_y[2904] = c_Body_y[2903];
                    end else begin
                        n_Body_x[2904] = c_Body_x[c_Size-1];
                        n_Body_y[2904] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2905) begin
                        n_Body_x[2905] = c_Body_x[2904];
                        n_Body_y[2905] = c_Body_y[2904];
                    end else begin
                        n_Body_x[2905] = c_Body_x[c_Size-1];
                        n_Body_y[2905] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2906) begin
                        n_Body_x[2906] = c_Body_x[2905];
                        n_Body_y[2906] = c_Body_y[2905];
                    end else begin
                        n_Body_x[2906] = c_Body_x[c_Size-1];
                        n_Body_y[2906] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2907) begin
                        n_Body_x[2907] = c_Body_x[2906];
                        n_Body_y[2907] = c_Body_y[2906];
                    end else begin
                        n_Body_x[2907] = c_Body_x[c_Size-1];
                        n_Body_y[2907] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2908) begin
                        n_Body_x[2908] = c_Body_x[2907];
                        n_Body_y[2908] = c_Body_y[2907];
                    end else begin
                        n_Body_x[2908] = c_Body_x[c_Size-1];
                        n_Body_y[2908] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2909) begin
                        n_Body_x[2909] = c_Body_x[2908];
                        n_Body_y[2909] = c_Body_y[2908];
                    end else begin
                        n_Body_x[2909] = c_Body_x[c_Size-1];
                        n_Body_y[2909] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2910) begin
                        n_Body_x[2910] = c_Body_x[2909];
                        n_Body_y[2910] = c_Body_y[2909];
                    end else begin
                        n_Body_x[2910] = c_Body_x[c_Size-1];
                        n_Body_y[2910] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2911) begin
                        n_Body_x[2911] = c_Body_x[2910];
                        n_Body_y[2911] = c_Body_y[2910];
                    end else begin
                        n_Body_x[2911] = c_Body_x[c_Size-1];
                        n_Body_y[2911] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2912) begin
                        n_Body_x[2912] = c_Body_x[2911];
                        n_Body_y[2912] = c_Body_y[2911];
                    end else begin
                        n_Body_x[2912] = c_Body_x[c_Size-1];
                        n_Body_y[2912] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2913) begin
                        n_Body_x[2913] = c_Body_x[2912];
                        n_Body_y[2913] = c_Body_y[2912];
                    end else begin
                        n_Body_x[2913] = c_Body_x[c_Size-1];
                        n_Body_y[2913] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2914) begin
                        n_Body_x[2914] = c_Body_x[2913];
                        n_Body_y[2914] = c_Body_y[2913];
                    end else begin
                        n_Body_x[2914] = c_Body_x[c_Size-1];
                        n_Body_y[2914] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2915) begin
                        n_Body_x[2915] = c_Body_x[2914];
                        n_Body_y[2915] = c_Body_y[2914];
                    end else begin
                        n_Body_x[2915] = c_Body_x[c_Size-1];
                        n_Body_y[2915] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2916) begin
                        n_Body_x[2916] = c_Body_x[2915];
                        n_Body_y[2916] = c_Body_y[2915];
                    end else begin
                        n_Body_x[2916] = c_Body_x[c_Size-1];
                        n_Body_y[2916] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2917) begin
                        n_Body_x[2917] = c_Body_x[2916];
                        n_Body_y[2917] = c_Body_y[2916];
                    end else begin
                        n_Body_x[2917] = c_Body_x[c_Size-1];
                        n_Body_y[2917] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2918) begin
                        n_Body_x[2918] = c_Body_x[2917];
                        n_Body_y[2918] = c_Body_y[2917];
                    end else begin
                        n_Body_x[2918] = c_Body_x[c_Size-1];
                        n_Body_y[2918] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2919) begin
                        n_Body_x[2919] = c_Body_x[2918];
                        n_Body_y[2919] = c_Body_y[2918];
                    end else begin
                        n_Body_x[2919] = c_Body_x[c_Size-1];
                        n_Body_y[2919] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2920) begin
                        n_Body_x[2920] = c_Body_x[2919];
                        n_Body_y[2920] = c_Body_y[2919];
                    end else begin
                        n_Body_x[2920] = c_Body_x[c_Size-1];
                        n_Body_y[2920] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2921) begin
                        n_Body_x[2921] = c_Body_x[2920];
                        n_Body_y[2921] = c_Body_y[2920];
                    end else begin
                        n_Body_x[2921] = c_Body_x[c_Size-1];
                        n_Body_y[2921] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2922) begin
                        n_Body_x[2922] = c_Body_x[2921];
                        n_Body_y[2922] = c_Body_y[2921];
                    end else begin
                        n_Body_x[2922] = c_Body_x[c_Size-1];
                        n_Body_y[2922] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2923) begin
                        n_Body_x[2923] = c_Body_x[2922];
                        n_Body_y[2923] = c_Body_y[2922];
                    end else begin
                        n_Body_x[2923] = c_Body_x[c_Size-1];
                        n_Body_y[2923] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2924) begin
                        n_Body_x[2924] = c_Body_x[2923];
                        n_Body_y[2924] = c_Body_y[2923];
                    end else begin
                        n_Body_x[2924] = c_Body_x[c_Size-1];
                        n_Body_y[2924] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2925) begin
                        n_Body_x[2925] = c_Body_x[2924];
                        n_Body_y[2925] = c_Body_y[2924];
                    end else begin
                        n_Body_x[2925] = c_Body_x[c_Size-1];
                        n_Body_y[2925] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2926) begin
                        n_Body_x[2926] = c_Body_x[2925];
                        n_Body_y[2926] = c_Body_y[2925];
                    end else begin
                        n_Body_x[2926] = c_Body_x[c_Size-1];
                        n_Body_y[2926] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2927) begin
                        n_Body_x[2927] = c_Body_x[2926];
                        n_Body_y[2927] = c_Body_y[2926];
                    end else begin
                        n_Body_x[2927] = c_Body_x[c_Size-1];
                        n_Body_y[2927] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2928) begin
                        n_Body_x[2928] = c_Body_x[2927];
                        n_Body_y[2928] = c_Body_y[2927];
                    end else begin
                        n_Body_x[2928] = c_Body_x[c_Size-1];
                        n_Body_y[2928] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2929) begin
                        n_Body_x[2929] = c_Body_x[2928];
                        n_Body_y[2929] = c_Body_y[2928];
                    end else begin
                        n_Body_x[2929] = c_Body_x[c_Size-1];
                        n_Body_y[2929] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2930) begin
                        n_Body_x[2930] = c_Body_x[2929];
                        n_Body_y[2930] = c_Body_y[2929];
                    end else begin
                        n_Body_x[2930] = c_Body_x[c_Size-1];
                        n_Body_y[2930] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2931) begin
                        n_Body_x[2931] = c_Body_x[2930];
                        n_Body_y[2931] = c_Body_y[2930];
                    end else begin
                        n_Body_x[2931] = c_Body_x[c_Size-1];
                        n_Body_y[2931] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2932) begin
                        n_Body_x[2932] = c_Body_x[2931];
                        n_Body_y[2932] = c_Body_y[2931];
                    end else begin
                        n_Body_x[2932] = c_Body_x[c_Size-1];
                        n_Body_y[2932] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2933) begin
                        n_Body_x[2933] = c_Body_x[2932];
                        n_Body_y[2933] = c_Body_y[2932];
                    end else begin
                        n_Body_x[2933] = c_Body_x[c_Size-1];
                        n_Body_y[2933] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2934) begin
                        n_Body_x[2934] = c_Body_x[2933];
                        n_Body_y[2934] = c_Body_y[2933];
                    end else begin
                        n_Body_x[2934] = c_Body_x[c_Size-1];
                        n_Body_y[2934] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2935) begin
                        n_Body_x[2935] = c_Body_x[2934];
                        n_Body_y[2935] = c_Body_y[2934];
                    end else begin
                        n_Body_x[2935] = c_Body_x[c_Size-1];
                        n_Body_y[2935] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2936) begin
                        n_Body_x[2936] = c_Body_x[2935];
                        n_Body_y[2936] = c_Body_y[2935];
                    end else begin
                        n_Body_x[2936] = c_Body_x[c_Size-1];
                        n_Body_y[2936] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2937) begin
                        n_Body_x[2937] = c_Body_x[2936];
                        n_Body_y[2937] = c_Body_y[2936];
                    end else begin
                        n_Body_x[2937] = c_Body_x[c_Size-1];
                        n_Body_y[2937] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2938) begin
                        n_Body_x[2938] = c_Body_x[2937];
                        n_Body_y[2938] = c_Body_y[2937];
                    end else begin
                        n_Body_x[2938] = c_Body_x[c_Size-1];
                        n_Body_y[2938] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2939) begin
                        n_Body_x[2939] = c_Body_x[2938];
                        n_Body_y[2939] = c_Body_y[2938];
                    end else begin
                        n_Body_x[2939] = c_Body_x[c_Size-1];
                        n_Body_y[2939] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2940) begin
                        n_Body_x[2940] = c_Body_x[2939];
                        n_Body_y[2940] = c_Body_y[2939];
                    end else begin
                        n_Body_x[2940] = c_Body_x[c_Size-1];
                        n_Body_y[2940] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2941) begin
                        n_Body_x[2941] = c_Body_x[2940];
                        n_Body_y[2941] = c_Body_y[2940];
                    end else begin
                        n_Body_x[2941] = c_Body_x[c_Size-1];
                        n_Body_y[2941] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2942) begin
                        n_Body_x[2942] = c_Body_x[2941];
                        n_Body_y[2942] = c_Body_y[2941];
                    end else begin
                        n_Body_x[2942] = c_Body_x[c_Size-1];
                        n_Body_y[2942] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2943) begin
                        n_Body_x[2943] = c_Body_x[2942];
                        n_Body_y[2943] = c_Body_y[2942];
                    end else begin
                        n_Body_x[2943] = c_Body_x[c_Size-1];
                        n_Body_y[2943] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2944) begin
                        n_Body_x[2944] = c_Body_x[2943];
                        n_Body_y[2944] = c_Body_y[2943];
                    end else begin
                        n_Body_x[2944] = c_Body_x[c_Size-1];
                        n_Body_y[2944] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2945) begin
                        n_Body_x[2945] = c_Body_x[2944];
                        n_Body_y[2945] = c_Body_y[2944];
                    end else begin
                        n_Body_x[2945] = c_Body_x[c_Size-1];
                        n_Body_y[2945] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2946) begin
                        n_Body_x[2946] = c_Body_x[2945];
                        n_Body_y[2946] = c_Body_y[2945];
                    end else begin
                        n_Body_x[2946] = c_Body_x[c_Size-1];
                        n_Body_y[2946] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2947) begin
                        n_Body_x[2947] = c_Body_x[2946];
                        n_Body_y[2947] = c_Body_y[2946];
                    end else begin
                        n_Body_x[2947] = c_Body_x[c_Size-1];
                        n_Body_y[2947] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2948) begin
                        n_Body_x[2948] = c_Body_x[2947];
                        n_Body_y[2948] = c_Body_y[2947];
                    end else begin
                        n_Body_x[2948] = c_Body_x[c_Size-1];
                        n_Body_y[2948] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2949) begin
                        n_Body_x[2949] = c_Body_x[2948];
                        n_Body_y[2949] = c_Body_y[2948];
                    end else begin
                        n_Body_x[2949] = c_Body_x[c_Size-1];
                        n_Body_y[2949] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2950) begin
                        n_Body_x[2950] = c_Body_x[2949];
                        n_Body_y[2950] = c_Body_y[2949];
                    end else begin
                        n_Body_x[2950] = c_Body_x[c_Size-1];
                        n_Body_y[2950] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2951) begin
                        n_Body_x[2951] = c_Body_x[2950];
                        n_Body_y[2951] = c_Body_y[2950];
                    end else begin
                        n_Body_x[2951] = c_Body_x[c_Size-1];
                        n_Body_y[2951] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2952) begin
                        n_Body_x[2952] = c_Body_x[2951];
                        n_Body_y[2952] = c_Body_y[2951];
                    end else begin
                        n_Body_x[2952] = c_Body_x[c_Size-1];
                        n_Body_y[2952] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2953) begin
                        n_Body_x[2953] = c_Body_x[2952];
                        n_Body_y[2953] = c_Body_y[2952];
                    end else begin
                        n_Body_x[2953] = c_Body_x[c_Size-1];
                        n_Body_y[2953] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2954) begin
                        n_Body_x[2954] = c_Body_x[2953];
                        n_Body_y[2954] = c_Body_y[2953];
                    end else begin
                        n_Body_x[2954] = c_Body_x[c_Size-1];
                        n_Body_y[2954] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2955) begin
                        n_Body_x[2955] = c_Body_x[2954];
                        n_Body_y[2955] = c_Body_y[2954];
                    end else begin
                        n_Body_x[2955] = c_Body_x[c_Size-1];
                        n_Body_y[2955] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2956) begin
                        n_Body_x[2956] = c_Body_x[2955];
                        n_Body_y[2956] = c_Body_y[2955];
                    end else begin
                        n_Body_x[2956] = c_Body_x[c_Size-1];
                        n_Body_y[2956] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2957) begin
                        n_Body_x[2957] = c_Body_x[2956];
                        n_Body_y[2957] = c_Body_y[2956];
                    end else begin
                        n_Body_x[2957] = c_Body_x[c_Size-1];
                        n_Body_y[2957] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2958) begin
                        n_Body_x[2958] = c_Body_x[2957];
                        n_Body_y[2958] = c_Body_y[2957];
                    end else begin
                        n_Body_x[2958] = c_Body_x[c_Size-1];
                        n_Body_y[2958] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2959) begin
                        n_Body_x[2959] = c_Body_x[2958];
                        n_Body_y[2959] = c_Body_y[2958];
                    end else begin
                        n_Body_x[2959] = c_Body_x[c_Size-1];
                        n_Body_y[2959] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2960) begin
                        n_Body_x[2960] = c_Body_x[2959];
                        n_Body_y[2960] = c_Body_y[2959];
                    end else begin
                        n_Body_x[2960] = c_Body_x[c_Size-1];
                        n_Body_y[2960] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2961) begin
                        n_Body_x[2961] = c_Body_x[2960];
                        n_Body_y[2961] = c_Body_y[2960];
                    end else begin
                        n_Body_x[2961] = c_Body_x[c_Size-1];
                        n_Body_y[2961] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2962) begin
                        n_Body_x[2962] = c_Body_x[2961];
                        n_Body_y[2962] = c_Body_y[2961];
                    end else begin
                        n_Body_x[2962] = c_Body_x[c_Size-1];
                        n_Body_y[2962] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2963) begin
                        n_Body_x[2963] = c_Body_x[2962];
                        n_Body_y[2963] = c_Body_y[2962];
                    end else begin
                        n_Body_x[2963] = c_Body_x[c_Size-1];
                        n_Body_y[2963] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2964) begin
                        n_Body_x[2964] = c_Body_x[2963];
                        n_Body_y[2964] = c_Body_y[2963];
                    end else begin
                        n_Body_x[2964] = c_Body_x[c_Size-1];
                        n_Body_y[2964] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2965) begin
                        n_Body_x[2965] = c_Body_x[2964];
                        n_Body_y[2965] = c_Body_y[2964];
                    end else begin
                        n_Body_x[2965] = c_Body_x[c_Size-1];
                        n_Body_y[2965] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2966) begin
                        n_Body_x[2966] = c_Body_x[2965];
                        n_Body_y[2966] = c_Body_y[2965];
                    end else begin
                        n_Body_x[2966] = c_Body_x[c_Size-1];
                        n_Body_y[2966] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2967) begin
                        n_Body_x[2967] = c_Body_x[2966];
                        n_Body_y[2967] = c_Body_y[2966];
                    end else begin
                        n_Body_x[2967] = c_Body_x[c_Size-1];
                        n_Body_y[2967] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2968) begin
                        n_Body_x[2968] = c_Body_x[2967];
                        n_Body_y[2968] = c_Body_y[2967];
                    end else begin
                        n_Body_x[2968] = c_Body_x[c_Size-1];
                        n_Body_y[2968] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2969) begin
                        n_Body_x[2969] = c_Body_x[2968];
                        n_Body_y[2969] = c_Body_y[2968];
                    end else begin
                        n_Body_x[2969] = c_Body_x[c_Size-1];
                        n_Body_y[2969] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2970) begin
                        n_Body_x[2970] = c_Body_x[2969];
                        n_Body_y[2970] = c_Body_y[2969];
                    end else begin
                        n_Body_x[2970] = c_Body_x[c_Size-1];
                        n_Body_y[2970] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2971) begin
                        n_Body_x[2971] = c_Body_x[2970];
                        n_Body_y[2971] = c_Body_y[2970];
                    end else begin
                        n_Body_x[2971] = c_Body_x[c_Size-1];
                        n_Body_y[2971] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2972) begin
                        n_Body_x[2972] = c_Body_x[2971];
                        n_Body_y[2972] = c_Body_y[2971];
                    end else begin
                        n_Body_x[2972] = c_Body_x[c_Size-1];
                        n_Body_y[2972] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2973) begin
                        n_Body_x[2973] = c_Body_x[2972];
                        n_Body_y[2973] = c_Body_y[2972];
                    end else begin
                        n_Body_x[2973] = c_Body_x[c_Size-1];
                        n_Body_y[2973] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2974) begin
                        n_Body_x[2974] = c_Body_x[2973];
                        n_Body_y[2974] = c_Body_y[2973];
                    end else begin
                        n_Body_x[2974] = c_Body_x[c_Size-1];
                        n_Body_y[2974] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2975) begin
                        n_Body_x[2975] = c_Body_x[2974];
                        n_Body_y[2975] = c_Body_y[2974];
                    end else begin
                        n_Body_x[2975] = c_Body_x[c_Size-1];
                        n_Body_y[2975] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2976) begin
                        n_Body_x[2976] = c_Body_x[2975];
                        n_Body_y[2976] = c_Body_y[2975];
                    end else begin
                        n_Body_x[2976] = c_Body_x[c_Size-1];
                        n_Body_y[2976] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2977) begin
                        n_Body_x[2977] = c_Body_x[2976];
                        n_Body_y[2977] = c_Body_y[2976];
                    end else begin
                        n_Body_x[2977] = c_Body_x[c_Size-1];
                        n_Body_y[2977] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2978) begin
                        n_Body_x[2978] = c_Body_x[2977];
                        n_Body_y[2978] = c_Body_y[2977];
                    end else begin
                        n_Body_x[2978] = c_Body_x[c_Size-1];
                        n_Body_y[2978] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2979) begin
                        n_Body_x[2979] = c_Body_x[2978];
                        n_Body_y[2979] = c_Body_y[2978];
                    end else begin
                        n_Body_x[2979] = c_Body_x[c_Size-1];
                        n_Body_y[2979] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2980) begin
                        n_Body_x[2980] = c_Body_x[2979];
                        n_Body_y[2980] = c_Body_y[2979];
                    end else begin
                        n_Body_x[2980] = c_Body_x[c_Size-1];
                        n_Body_y[2980] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2981) begin
                        n_Body_x[2981] = c_Body_x[2980];
                        n_Body_y[2981] = c_Body_y[2980];
                    end else begin
                        n_Body_x[2981] = c_Body_x[c_Size-1];
                        n_Body_y[2981] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2982) begin
                        n_Body_x[2982] = c_Body_x[2981];
                        n_Body_y[2982] = c_Body_y[2981];
                    end else begin
                        n_Body_x[2982] = c_Body_x[c_Size-1];
                        n_Body_y[2982] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2983) begin
                        n_Body_x[2983] = c_Body_x[2982];
                        n_Body_y[2983] = c_Body_y[2982];
                    end else begin
                        n_Body_x[2983] = c_Body_x[c_Size-1];
                        n_Body_y[2983] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2984) begin
                        n_Body_x[2984] = c_Body_x[2983];
                        n_Body_y[2984] = c_Body_y[2983];
                    end else begin
                        n_Body_x[2984] = c_Body_x[c_Size-1];
                        n_Body_y[2984] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2985) begin
                        n_Body_x[2985] = c_Body_x[2984];
                        n_Body_y[2985] = c_Body_y[2984];
                    end else begin
                        n_Body_x[2985] = c_Body_x[c_Size-1];
                        n_Body_y[2985] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2986) begin
                        n_Body_x[2986] = c_Body_x[2985];
                        n_Body_y[2986] = c_Body_y[2985];
                    end else begin
                        n_Body_x[2986] = c_Body_x[c_Size-1];
                        n_Body_y[2986] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2987) begin
                        n_Body_x[2987] = c_Body_x[2986];
                        n_Body_y[2987] = c_Body_y[2986];
                    end else begin
                        n_Body_x[2987] = c_Body_x[c_Size-1];
                        n_Body_y[2987] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2988) begin
                        n_Body_x[2988] = c_Body_x[2987];
                        n_Body_y[2988] = c_Body_y[2987];
                    end else begin
                        n_Body_x[2988] = c_Body_x[c_Size-1];
                        n_Body_y[2988] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2989) begin
                        n_Body_x[2989] = c_Body_x[2988];
                        n_Body_y[2989] = c_Body_y[2988];
                    end else begin
                        n_Body_x[2989] = c_Body_x[c_Size-1];
                        n_Body_y[2989] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2990) begin
                        n_Body_x[2990] = c_Body_x[2989];
                        n_Body_y[2990] = c_Body_y[2989];
                    end else begin
                        n_Body_x[2990] = c_Body_x[c_Size-1];
                        n_Body_y[2990] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2991) begin
                        n_Body_x[2991] = c_Body_x[2990];
                        n_Body_y[2991] = c_Body_y[2990];
                    end else begin
                        n_Body_x[2991] = c_Body_x[c_Size-1];
                        n_Body_y[2991] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2992) begin
                        n_Body_x[2992] = c_Body_x[2991];
                        n_Body_y[2992] = c_Body_y[2991];
                    end else begin
                        n_Body_x[2992] = c_Body_x[c_Size-1];
                        n_Body_y[2992] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2993) begin
                        n_Body_x[2993] = c_Body_x[2992];
                        n_Body_y[2993] = c_Body_y[2992];
                    end else begin
                        n_Body_x[2993] = c_Body_x[c_Size-1];
                        n_Body_y[2993] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2994) begin
                        n_Body_x[2994] = c_Body_x[2993];
                        n_Body_y[2994] = c_Body_y[2993];
                    end else begin
                        n_Body_x[2994] = c_Body_x[c_Size-1];
                        n_Body_y[2994] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2995) begin
                        n_Body_x[2995] = c_Body_x[2994];
                        n_Body_y[2995] = c_Body_y[2994];
                    end else begin
                        n_Body_x[2995] = c_Body_x[c_Size-1];
                        n_Body_y[2995] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2996) begin
                        n_Body_x[2996] = c_Body_x[2995];
                        n_Body_y[2996] = c_Body_y[2995];
                    end else begin
                        n_Body_x[2996] = c_Body_x[c_Size-1];
                        n_Body_y[2996] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2997) begin
                        n_Body_x[2997] = c_Body_x[2996];
                        n_Body_y[2997] = c_Body_y[2996];
                    end else begin
                        n_Body_x[2997] = c_Body_x[c_Size-1];
                        n_Body_y[2997] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2998) begin
                        n_Body_x[2998] = c_Body_x[2997];
                        n_Body_y[2998] = c_Body_y[2997];
                    end else begin
                        n_Body_x[2998] = c_Body_x[c_Size-1];
                        n_Body_y[2998] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 2999) begin
                        n_Body_x[2999] = c_Body_x[2998];
                        n_Body_y[2999] = c_Body_y[2998];
                    end else begin
                        n_Body_x[2999] = c_Body_x[c_Size-1];
                        n_Body_y[2999] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3000) begin
                        n_Body_x[3000] = c_Body_x[2999];
                        n_Body_y[3000] = c_Body_y[2999];
                    end else begin
                        n_Body_x[3000] = c_Body_x[c_Size-1];
                        n_Body_y[3000] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3001) begin
                        n_Body_x[3001] = c_Body_x[3000];
                        n_Body_y[3001] = c_Body_y[3000];
                    end else begin
                        n_Body_x[3001] = c_Body_x[c_Size-1];
                        n_Body_y[3001] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3002) begin
                        n_Body_x[3002] = c_Body_x[3001];
                        n_Body_y[3002] = c_Body_y[3001];
                    end else begin
                        n_Body_x[3002] = c_Body_x[c_Size-1];
                        n_Body_y[3002] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3003) begin
                        n_Body_x[3003] = c_Body_x[3002];
                        n_Body_y[3003] = c_Body_y[3002];
                    end else begin
                        n_Body_x[3003] = c_Body_x[c_Size-1];
                        n_Body_y[3003] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3004) begin
                        n_Body_x[3004] = c_Body_x[3003];
                        n_Body_y[3004] = c_Body_y[3003];
                    end else begin
                        n_Body_x[3004] = c_Body_x[c_Size-1];
                        n_Body_y[3004] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3005) begin
                        n_Body_x[3005] = c_Body_x[3004];
                        n_Body_y[3005] = c_Body_y[3004];
                    end else begin
                        n_Body_x[3005] = c_Body_x[c_Size-1];
                        n_Body_y[3005] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3006) begin
                        n_Body_x[3006] = c_Body_x[3005];
                        n_Body_y[3006] = c_Body_y[3005];
                    end else begin
                        n_Body_x[3006] = c_Body_x[c_Size-1];
                        n_Body_y[3006] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3007) begin
                        n_Body_x[3007] = c_Body_x[3006];
                        n_Body_y[3007] = c_Body_y[3006];
                    end else begin
                        n_Body_x[3007] = c_Body_x[c_Size-1];
                        n_Body_y[3007] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3008) begin
                        n_Body_x[3008] = c_Body_x[3007];
                        n_Body_y[3008] = c_Body_y[3007];
                    end else begin
                        n_Body_x[3008] = c_Body_x[c_Size-1];
                        n_Body_y[3008] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3009) begin
                        n_Body_x[3009] = c_Body_x[3008];
                        n_Body_y[3009] = c_Body_y[3008];
                    end else begin
                        n_Body_x[3009] = c_Body_x[c_Size-1];
                        n_Body_y[3009] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3010) begin
                        n_Body_x[3010] = c_Body_x[3009];
                        n_Body_y[3010] = c_Body_y[3009];
                    end else begin
                        n_Body_x[3010] = c_Body_x[c_Size-1];
                        n_Body_y[3010] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3011) begin
                        n_Body_x[3011] = c_Body_x[3010];
                        n_Body_y[3011] = c_Body_y[3010];
                    end else begin
                        n_Body_x[3011] = c_Body_x[c_Size-1];
                        n_Body_y[3011] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3012) begin
                        n_Body_x[3012] = c_Body_x[3011];
                        n_Body_y[3012] = c_Body_y[3011];
                    end else begin
                        n_Body_x[3012] = c_Body_x[c_Size-1];
                        n_Body_y[3012] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3013) begin
                        n_Body_x[3013] = c_Body_x[3012];
                        n_Body_y[3013] = c_Body_y[3012];
                    end else begin
                        n_Body_x[3013] = c_Body_x[c_Size-1];
                        n_Body_y[3013] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3014) begin
                        n_Body_x[3014] = c_Body_x[3013];
                        n_Body_y[3014] = c_Body_y[3013];
                    end else begin
                        n_Body_x[3014] = c_Body_x[c_Size-1];
                        n_Body_y[3014] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3015) begin
                        n_Body_x[3015] = c_Body_x[3014];
                        n_Body_y[3015] = c_Body_y[3014];
                    end else begin
                        n_Body_x[3015] = c_Body_x[c_Size-1];
                        n_Body_y[3015] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3016) begin
                        n_Body_x[3016] = c_Body_x[3015];
                        n_Body_y[3016] = c_Body_y[3015];
                    end else begin
                        n_Body_x[3016] = c_Body_x[c_Size-1];
                        n_Body_y[3016] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3017) begin
                        n_Body_x[3017] = c_Body_x[3016];
                        n_Body_y[3017] = c_Body_y[3016];
                    end else begin
                        n_Body_x[3017] = c_Body_x[c_Size-1];
                        n_Body_y[3017] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3018) begin
                        n_Body_x[3018] = c_Body_x[3017];
                        n_Body_y[3018] = c_Body_y[3017];
                    end else begin
                        n_Body_x[3018] = c_Body_x[c_Size-1];
                        n_Body_y[3018] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3019) begin
                        n_Body_x[3019] = c_Body_x[3018];
                        n_Body_y[3019] = c_Body_y[3018];
                    end else begin
                        n_Body_x[3019] = c_Body_x[c_Size-1];
                        n_Body_y[3019] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3020) begin
                        n_Body_x[3020] = c_Body_x[3019];
                        n_Body_y[3020] = c_Body_y[3019];
                    end else begin
                        n_Body_x[3020] = c_Body_x[c_Size-1];
                        n_Body_y[3020] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3021) begin
                        n_Body_x[3021] = c_Body_x[3020];
                        n_Body_y[3021] = c_Body_y[3020];
                    end else begin
                        n_Body_x[3021] = c_Body_x[c_Size-1];
                        n_Body_y[3021] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3022) begin
                        n_Body_x[3022] = c_Body_x[3021];
                        n_Body_y[3022] = c_Body_y[3021];
                    end else begin
                        n_Body_x[3022] = c_Body_x[c_Size-1];
                        n_Body_y[3022] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3023) begin
                        n_Body_x[3023] = c_Body_x[3022];
                        n_Body_y[3023] = c_Body_y[3022];
                    end else begin
                        n_Body_x[3023] = c_Body_x[c_Size-1];
                        n_Body_y[3023] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3024) begin
                        n_Body_x[3024] = c_Body_x[3023];
                        n_Body_y[3024] = c_Body_y[3023];
                    end else begin
                        n_Body_x[3024] = c_Body_x[c_Size-1];
                        n_Body_y[3024] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3025) begin
                        n_Body_x[3025] = c_Body_x[3024];
                        n_Body_y[3025] = c_Body_y[3024];
                    end else begin
                        n_Body_x[3025] = c_Body_x[c_Size-1];
                        n_Body_y[3025] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3026) begin
                        n_Body_x[3026] = c_Body_x[3025];
                        n_Body_y[3026] = c_Body_y[3025];
                    end else begin
                        n_Body_x[3026] = c_Body_x[c_Size-1];
                        n_Body_y[3026] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3027) begin
                        n_Body_x[3027] = c_Body_x[3026];
                        n_Body_y[3027] = c_Body_y[3026];
                    end else begin
                        n_Body_x[3027] = c_Body_x[c_Size-1];
                        n_Body_y[3027] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3028) begin
                        n_Body_x[3028] = c_Body_x[3027];
                        n_Body_y[3028] = c_Body_y[3027];
                    end else begin
                        n_Body_x[3028] = c_Body_x[c_Size-1];
                        n_Body_y[3028] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3029) begin
                        n_Body_x[3029] = c_Body_x[3028];
                        n_Body_y[3029] = c_Body_y[3028];
                    end else begin
                        n_Body_x[3029] = c_Body_x[c_Size-1];
                        n_Body_y[3029] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3030) begin
                        n_Body_x[3030] = c_Body_x[3029];
                        n_Body_y[3030] = c_Body_y[3029];
                    end else begin
                        n_Body_x[3030] = c_Body_x[c_Size-1];
                        n_Body_y[3030] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3031) begin
                        n_Body_x[3031] = c_Body_x[3030];
                        n_Body_y[3031] = c_Body_y[3030];
                    end else begin
                        n_Body_x[3031] = c_Body_x[c_Size-1];
                        n_Body_y[3031] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3032) begin
                        n_Body_x[3032] = c_Body_x[3031];
                        n_Body_y[3032] = c_Body_y[3031];
                    end else begin
                        n_Body_x[3032] = c_Body_x[c_Size-1];
                        n_Body_y[3032] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3033) begin
                        n_Body_x[3033] = c_Body_x[3032];
                        n_Body_y[3033] = c_Body_y[3032];
                    end else begin
                        n_Body_x[3033] = c_Body_x[c_Size-1];
                        n_Body_y[3033] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3034) begin
                        n_Body_x[3034] = c_Body_x[3033];
                        n_Body_y[3034] = c_Body_y[3033];
                    end else begin
                        n_Body_x[3034] = c_Body_x[c_Size-1];
                        n_Body_y[3034] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3035) begin
                        n_Body_x[3035] = c_Body_x[3034];
                        n_Body_y[3035] = c_Body_y[3034];
                    end else begin
                        n_Body_x[3035] = c_Body_x[c_Size-1];
                        n_Body_y[3035] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3036) begin
                        n_Body_x[3036] = c_Body_x[3035];
                        n_Body_y[3036] = c_Body_y[3035];
                    end else begin
                        n_Body_x[3036] = c_Body_x[c_Size-1];
                        n_Body_y[3036] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3037) begin
                        n_Body_x[3037] = c_Body_x[3036];
                        n_Body_y[3037] = c_Body_y[3036];
                    end else begin
                        n_Body_x[3037] = c_Body_x[c_Size-1];
                        n_Body_y[3037] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3038) begin
                        n_Body_x[3038] = c_Body_x[3037];
                        n_Body_y[3038] = c_Body_y[3037];
                    end else begin
                        n_Body_x[3038] = c_Body_x[c_Size-1];
                        n_Body_y[3038] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3039) begin
                        n_Body_x[3039] = c_Body_x[3038];
                        n_Body_y[3039] = c_Body_y[3038];
                    end else begin
                        n_Body_x[3039] = c_Body_x[c_Size-1];
                        n_Body_y[3039] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3040) begin
                        n_Body_x[3040] = c_Body_x[3039];
                        n_Body_y[3040] = c_Body_y[3039];
                    end else begin
                        n_Body_x[3040] = c_Body_x[c_Size-1];
                        n_Body_y[3040] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3041) begin
                        n_Body_x[3041] = c_Body_x[3040];
                        n_Body_y[3041] = c_Body_y[3040];
                    end else begin
                        n_Body_x[3041] = c_Body_x[c_Size-1];
                        n_Body_y[3041] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3042) begin
                        n_Body_x[3042] = c_Body_x[3041];
                        n_Body_y[3042] = c_Body_y[3041];
                    end else begin
                        n_Body_x[3042] = c_Body_x[c_Size-1];
                        n_Body_y[3042] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3043) begin
                        n_Body_x[3043] = c_Body_x[3042];
                        n_Body_y[3043] = c_Body_y[3042];
                    end else begin
                        n_Body_x[3043] = c_Body_x[c_Size-1];
                        n_Body_y[3043] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3044) begin
                        n_Body_x[3044] = c_Body_x[3043];
                        n_Body_y[3044] = c_Body_y[3043];
                    end else begin
                        n_Body_x[3044] = c_Body_x[c_Size-1];
                        n_Body_y[3044] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3045) begin
                        n_Body_x[3045] = c_Body_x[3044];
                        n_Body_y[3045] = c_Body_y[3044];
                    end else begin
                        n_Body_x[3045] = c_Body_x[c_Size-1];
                        n_Body_y[3045] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3046) begin
                        n_Body_x[3046] = c_Body_x[3045];
                        n_Body_y[3046] = c_Body_y[3045];
                    end else begin
                        n_Body_x[3046] = c_Body_x[c_Size-1];
                        n_Body_y[3046] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3047) begin
                        n_Body_x[3047] = c_Body_x[3046];
                        n_Body_y[3047] = c_Body_y[3046];
                    end else begin
                        n_Body_x[3047] = c_Body_x[c_Size-1];
                        n_Body_y[3047] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3048) begin
                        n_Body_x[3048] = c_Body_x[3047];
                        n_Body_y[3048] = c_Body_y[3047];
                    end else begin
                        n_Body_x[3048] = c_Body_x[c_Size-1];
                        n_Body_y[3048] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3049) begin
                        n_Body_x[3049] = c_Body_x[3048];
                        n_Body_y[3049] = c_Body_y[3048];
                    end else begin
                        n_Body_x[3049] = c_Body_x[c_Size-1];
                        n_Body_y[3049] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3050) begin
                        n_Body_x[3050] = c_Body_x[3049];
                        n_Body_y[3050] = c_Body_y[3049];
                    end else begin
                        n_Body_x[3050] = c_Body_x[c_Size-1];
                        n_Body_y[3050] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3051) begin
                        n_Body_x[3051] = c_Body_x[3050];
                        n_Body_y[3051] = c_Body_y[3050];
                    end else begin
                        n_Body_x[3051] = c_Body_x[c_Size-1];
                        n_Body_y[3051] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3052) begin
                        n_Body_x[3052] = c_Body_x[3051];
                        n_Body_y[3052] = c_Body_y[3051];
                    end else begin
                        n_Body_x[3052] = c_Body_x[c_Size-1];
                        n_Body_y[3052] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3053) begin
                        n_Body_x[3053] = c_Body_x[3052];
                        n_Body_y[3053] = c_Body_y[3052];
                    end else begin
                        n_Body_x[3053] = c_Body_x[c_Size-1];
                        n_Body_y[3053] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3054) begin
                        n_Body_x[3054] = c_Body_x[3053];
                        n_Body_y[3054] = c_Body_y[3053];
                    end else begin
                        n_Body_x[3054] = c_Body_x[c_Size-1];
                        n_Body_y[3054] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3055) begin
                        n_Body_x[3055] = c_Body_x[3054];
                        n_Body_y[3055] = c_Body_y[3054];
                    end else begin
                        n_Body_x[3055] = c_Body_x[c_Size-1];
                        n_Body_y[3055] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3056) begin
                        n_Body_x[3056] = c_Body_x[3055];
                        n_Body_y[3056] = c_Body_y[3055];
                    end else begin
                        n_Body_x[3056] = c_Body_x[c_Size-1];
                        n_Body_y[3056] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3057) begin
                        n_Body_x[3057] = c_Body_x[3056];
                        n_Body_y[3057] = c_Body_y[3056];
                    end else begin
                        n_Body_x[3057] = c_Body_x[c_Size-1];
                        n_Body_y[3057] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3058) begin
                        n_Body_x[3058] = c_Body_x[3057];
                        n_Body_y[3058] = c_Body_y[3057];
                    end else begin
                        n_Body_x[3058] = c_Body_x[c_Size-1];
                        n_Body_y[3058] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3059) begin
                        n_Body_x[3059] = c_Body_x[3058];
                        n_Body_y[3059] = c_Body_y[3058];
                    end else begin
                        n_Body_x[3059] = c_Body_x[c_Size-1];
                        n_Body_y[3059] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3060) begin
                        n_Body_x[3060] = c_Body_x[3059];
                        n_Body_y[3060] = c_Body_y[3059];
                    end else begin
                        n_Body_x[3060] = c_Body_x[c_Size-1];
                        n_Body_y[3060] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3061) begin
                        n_Body_x[3061] = c_Body_x[3060];
                        n_Body_y[3061] = c_Body_y[3060];
                    end else begin
                        n_Body_x[3061] = c_Body_x[c_Size-1];
                        n_Body_y[3061] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3062) begin
                        n_Body_x[3062] = c_Body_x[3061];
                        n_Body_y[3062] = c_Body_y[3061];
                    end else begin
                        n_Body_x[3062] = c_Body_x[c_Size-1];
                        n_Body_y[3062] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3063) begin
                        n_Body_x[3063] = c_Body_x[3062];
                        n_Body_y[3063] = c_Body_y[3062];
                    end else begin
                        n_Body_x[3063] = c_Body_x[c_Size-1];
                        n_Body_y[3063] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3064) begin
                        n_Body_x[3064] = c_Body_x[3063];
                        n_Body_y[3064] = c_Body_y[3063];
                    end else begin
                        n_Body_x[3064] = c_Body_x[c_Size-1];
                        n_Body_y[3064] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3065) begin
                        n_Body_x[3065] = c_Body_x[3064];
                        n_Body_y[3065] = c_Body_y[3064];
                    end else begin
                        n_Body_x[3065] = c_Body_x[c_Size-1];
                        n_Body_y[3065] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3066) begin
                        n_Body_x[3066] = c_Body_x[3065];
                        n_Body_y[3066] = c_Body_y[3065];
                    end else begin
                        n_Body_x[3066] = c_Body_x[c_Size-1];
                        n_Body_y[3066] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3067) begin
                        n_Body_x[3067] = c_Body_x[3066];
                        n_Body_y[3067] = c_Body_y[3066];
                    end else begin
                        n_Body_x[3067] = c_Body_x[c_Size-1];
                        n_Body_y[3067] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3068) begin
                        n_Body_x[3068] = c_Body_x[3067];
                        n_Body_y[3068] = c_Body_y[3067];
                    end else begin
                        n_Body_x[3068] = c_Body_x[c_Size-1];
                        n_Body_y[3068] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3069) begin
                        n_Body_x[3069] = c_Body_x[3068];
                        n_Body_y[3069] = c_Body_y[3068];
                    end else begin
                        n_Body_x[3069] = c_Body_x[c_Size-1];
                        n_Body_y[3069] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3070) begin
                        n_Body_x[3070] = c_Body_x[3069];
                        n_Body_y[3070] = c_Body_y[3069];
                    end else begin
                        n_Body_x[3070] = c_Body_x[c_Size-1];
                        n_Body_y[3070] = c_Body_y[c_Size-1];
                    end
                    if (n_Size > 3071) begin
                        n_Body_x[3071] = c_Body_x[3070];
                        n_Body_y[3071] = c_Body_y[3070];
                    end else begin
                        n_Body_x[3071] = c_Body_x[c_Size-1];
                        n_Body_y[3071] = c_Body_y[c_Size-1];
                    end
            end
            PAUSE : begin
                n_State = !i_Pause ? RUN : c_State;
            end
            STOP : begin

            end
        endcase
    end
endmodule