module Vga (
    i_Clk,            // 50 MHz 입력 클럭
    i_Rst,            // 리셋 신호
    i_worm_x,           // 지렁이 x 위치 배열
    i_worm_y,           // 지렁이 y 위치 배열
    i_item_x,           // 아이템의 x 위치 (0~64)
    i_item_y,           // 아이템의 y 위치 (0~48)
    i_size,
    o_hsync,            // 수평 동기 신호
    o_vsync,            // 수직 동기 신호
    o_red,              // 빨강 색상 데이터
    o_green,            // 초록 색상 데이터
    o_blue              // 파랑 색상 데이터
);
    
    input i_Clk;
    input i_Rst;

    parameter MAX_SIZE   = 3072;
    input [MAX_SIZE * 6 - 1:0] i_worm_x;
    input [MAX_SIZE * 6 - 1:0] i_worm_y;

    input [5:0] i_item_x;
    input [5:0] i_item_y;

    input [11:0] i_size;

    output o_hsync;
    output o_vsync;

    output reg[7:0] o_red;
    output reg[7:0] o_green;
    output reg[7:0] o_blue;

    // 픽셀 클럭 분주 (50MHz -> 25MHz)
    reg pixel_clk;
    always @(posedge i_Clk or posedge i_Rst) begin
        if (i_Rst)
            pixel_clk <= 0;
        else
            pixel_clk <= ~pixel_clk;
    end

    // VGA 640x480 @ 60Hz (25.175 MHz 픽셀 클럭) 타이밍
    parameter H_DISPLAY = 640;
    parameter H_FRONT = 16;
    parameter H_SYNC = 96;
    parameter H_BACK = 48;
    parameter H_TOTAL = 800;

    parameter V_DISPLAY = 480;
    parameter V_FRONT = 10;
    parameter V_SYNC = 2;
    parameter V_BACK = 33;
    parameter V_TOTAL = 525;
    
    parameter PIXEL_SIZE = 10;

    reg [9:0] h_count; // 수평 픽셀 카운터
    reg [9:0] v_count; // 수직 픽셀 카운터
    reg worm_active;

    wire active_area = (h_count < H_DISPLAY) && (v_count < V_DISPLAY);

    // 동기 신호 생성
    assign o_hsync = ~(h_count >= (H_DISPLAY + H_FRONT) && h_count < (H_DISPLAY + H_FRONT + H_SYNC));
    assign o_vsync = ~(v_count >= (V_DISPLAY + V_FRONT) && v_count < (V_DISPLAY + V_FRONT + V_SYNC));

    // 아이템 위치 확대 스케일링
    wire [9:0] item_x_scaled = i_item_x * PIXEL_SIZE;
    wire [9:0] item_y_scaled = i_item_y * PIXEL_SIZE;

    wire item_active = h_count >= item_x_scaled && h_count < item_x_scaled + 10 &&
                       v_count >= item_y_scaled && v_count < item_y_scaled + 10;
    wire edge_active = h_count == 0 || h_count == H_DISPLAY - 1 ||
                       v_count == 0 || v_count == V_DISPLAY - 1;


    always @(posedge pixel_clk or posedge i_Rst) begin
        if (i_Rst) begin
            h_count = 0;
            v_count = 0;
            o_red = 0;
            o_green = 0;
            o_blue = 0;
            worm_active = 0;
        end else begin
            // 수평 및 수직 카운터
            if (h_count < H_TOTAL - 1) begin
                h_count = h_count + 1;
            end else begin
                h_count = 0;
                if (v_count < V_TOTAL - 1) begin
                    v_count = v_count + 1;
                end else begin
                    v_count = 0;
                end
            end

            // 픽셀 데이터 출력
            if (active_area) begin
                worm_active = 0;
                // 지렁이 배열 확인
                     if (0 < i_size && h_count >= i_worm_x[5:0] * PIXEL_SIZE && h_count < i_worm_x[5:0] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5:0] * PIXEL_SIZE && v_count < i_worm_y[5:0] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1 < i_size && h_count >= i_worm_x[11:6] * PIXEL_SIZE && h_count < i_worm_x[11:6] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11:6] * PIXEL_SIZE && v_count < i_worm_y[11:6] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2 < i_size && h_count >= i_worm_x[17:12] * PIXEL_SIZE && h_count < i_worm_x[17:12] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17:12] * PIXEL_SIZE && v_count < i_worm_y[17:12] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3 < i_size && h_count >= i_worm_x[23:18] * PIXEL_SIZE && h_count < i_worm_x[23:18] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[23:18] * PIXEL_SIZE && v_count < i_worm_y[23:18] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (4 < i_size && h_count >= i_worm_x[29:24] * PIXEL_SIZE && h_count < i_worm_x[29:24] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[29:24] * PIXEL_SIZE && v_count < i_worm_y[29:24] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (5 < i_size && h_count >= i_worm_x[35:30] * PIXEL_SIZE && h_count < i_worm_x[35:30] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[35:30] * PIXEL_SIZE && v_count < i_worm_y[35:30] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (6 < i_size && h_count >= i_worm_x[41:36] * PIXEL_SIZE && h_count < i_worm_x[41:36] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[41:36] * PIXEL_SIZE && v_count < i_worm_y[41:36] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (7 < i_size && h_count >= i_worm_x[47:42] * PIXEL_SIZE && h_count < i_worm_x[47:42] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[47:42] * PIXEL_SIZE && v_count < i_worm_y[47:42] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (8 < i_size && h_count >= i_worm_x[53:48] * PIXEL_SIZE && h_count < i_worm_x[53:48] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[53:48] * PIXEL_SIZE && v_count < i_worm_y[53:48] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (9 < i_size && h_count >= i_worm_x[59:54] * PIXEL_SIZE && h_count < i_worm_x[59:54] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[59:54] * PIXEL_SIZE && v_count < i_worm_y[59:54] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (10 < i_size && h_count >= i_worm_x[65:60] * PIXEL_SIZE && h_count < i_worm_x[65:60] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[65:60] * PIXEL_SIZE && v_count < i_worm_y[65:60] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (11 < i_size && h_count >= i_worm_x[71:66] * PIXEL_SIZE && h_count < i_worm_x[71:66] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[71:66] * PIXEL_SIZE && v_count < i_worm_y[71:66] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (12 < i_size && h_count >= i_worm_x[77:72] * PIXEL_SIZE && h_count < i_worm_x[77:72] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[77:72] * PIXEL_SIZE && v_count < i_worm_y[77:72] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (13 < i_size && h_count >= i_worm_x[83:78] * PIXEL_SIZE && h_count < i_worm_x[83:78] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[83:78] * PIXEL_SIZE && v_count < i_worm_y[83:78] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (14 < i_size && h_count >= i_worm_x[89:84] * PIXEL_SIZE && h_count < i_worm_x[89:84] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[89:84] * PIXEL_SIZE && v_count < i_worm_y[89:84] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (15 < i_size && h_count >= i_worm_x[95:90] * PIXEL_SIZE && h_count < i_worm_x[95:90] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[95:90] * PIXEL_SIZE && v_count < i_worm_y[95:90] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (16 < i_size && h_count >= i_worm_x[101:96] * PIXEL_SIZE && h_count < i_worm_x[101:96] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[101:96] * PIXEL_SIZE && v_count < i_worm_y[101:96] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (17 < i_size && h_count >= i_worm_x[107:102] * PIXEL_SIZE && h_count < i_worm_x[107:102] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[107:102] * PIXEL_SIZE && v_count < i_worm_y[107:102] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (18 < i_size && h_count >= i_worm_x[113:108] * PIXEL_SIZE && h_count < i_worm_x[113:108] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[113:108] * PIXEL_SIZE && v_count < i_worm_y[113:108] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (19 < i_size && h_count >= i_worm_x[119:114] * PIXEL_SIZE && h_count < i_worm_x[119:114] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[119:114] * PIXEL_SIZE && v_count < i_worm_y[119:114] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (20 < i_size && h_count >= i_worm_x[125:120] * PIXEL_SIZE && h_count < i_worm_x[125:120] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[125:120] * PIXEL_SIZE && v_count < i_worm_y[125:120] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (21 < i_size && h_count >= i_worm_x[131:126] * PIXEL_SIZE && h_count < i_worm_x[131:126] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[131:126] * PIXEL_SIZE && v_count < i_worm_y[131:126] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (22 < i_size && h_count >= i_worm_x[137:132] * PIXEL_SIZE && h_count < i_worm_x[137:132] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[137:132] * PIXEL_SIZE && v_count < i_worm_y[137:132] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (23 < i_size && h_count >= i_worm_x[143:138] * PIXEL_SIZE && h_count < i_worm_x[143:138] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[143:138] * PIXEL_SIZE && v_count < i_worm_y[143:138] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (24 < i_size && h_count >= i_worm_x[149:144] * PIXEL_SIZE && h_count < i_worm_x[149:144] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[149:144] * PIXEL_SIZE && v_count < i_worm_y[149:144] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (25 < i_size && h_count >= i_worm_x[155:150] * PIXEL_SIZE && h_count < i_worm_x[155:150] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[155:150] * PIXEL_SIZE && v_count < i_worm_y[155:150] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (26 < i_size && h_count >= i_worm_x[161:156] * PIXEL_SIZE && h_count < i_worm_x[161:156] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[161:156] * PIXEL_SIZE && v_count < i_worm_y[161:156] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (27 < i_size && h_count >= i_worm_x[167:162] * PIXEL_SIZE && h_count < i_worm_x[167:162] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[167:162] * PIXEL_SIZE && v_count < i_worm_y[167:162] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (28 < i_size && h_count >= i_worm_x[173:168] * PIXEL_SIZE && h_count < i_worm_x[173:168] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[173:168] * PIXEL_SIZE && v_count < i_worm_y[173:168] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (29 < i_size && h_count >= i_worm_x[179:174] * PIXEL_SIZE && h_count < i_worm_x[179:174] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[179:174] * PIXEL_SIZE && v_count < i_worm_y[179:174] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (30 < i_size && h_count >= i_worm_x[185:180] * PIXEL_SIZE && h_count < i_worm_x[185:180] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[185:180] * PIXEL_SIZE && v_count < i_worm_y[185:180] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (31 < i_size && h_count >= i_worm_x[191:186] * PIXEL_SIZE && h_count < i_worm_x[191:186] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[191:186] * PIXEL_SIZE && v_count < i_worm_y[191:186] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (32 < i_size && h_count >= i_worm_x[197:192] * PIXEL_SIZE && h_count < i_worm_x[197:192] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[197:192] * PIXEL_SIZE && v_count < i_worm_y[197:192] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (33 < i_size && h_count >= i_worm_x[203:198] * PIXEL_SIZE && h_count < i_worm_x[203:198] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[203:198] * PIXEL_SIZE && v_count < i_worm_y[203:198] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (34 < i_size && h_count >= i_worm_x[209:204] * PIXEL_SIZE && h_count < i_worm_x[209:204] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[209:204] * PIXEL_SIZE && v_count < i_worm_y[209:204] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (35 < i_size && h_count >= i_worm_x[215:210] * PIXEL_SIZE && h_count < i_worm_x[215:210] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[215:210] * PIXEL_SIZE && v_count < i_worm_y[215:210] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (36 < i_size && h_count >= i_worm_x[221:216] * PIXEL_SIZE && h_count < i_worm_x[221:216] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[221:216] * PIXEL_SIZE && v_count < i_worm_y[221:216] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (37 < i_size && h_count >= i_worm_x[227:222] * PIXEL_SIZE && h_count < i_worm_x[227:222] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[227:222] * PIXEL_SIZE && v_count < i_worm_y[227:222] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (38 < i_size && h_count >= i_worm_x[233:228] * PIXEL_SIZE && h_count < i_worm_x[233:228] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[233:228] * PIXEL_SIZE && v_count < i_worm_y[233:228] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (39 < i_size && h_count >= i_worm_x[239:234] * PIXEL_SIZE && h_count < i_worm_x[239:234] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[239:234] * PIXEL_SIZE && v_count < i_worm_y[239:234] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (40 < i_size && h_count >= i_worm_x[245:240] * PIXEL_SIZE && h_count < i_worm_x[245:240] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[245:240] * PIXEL_SIZE && v_count < i_worm_y[245:240] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (41 < i_size && h_count >= i_worm_x[251:246] * PIXEL_SIZE && h_count < i_worm_x[251:246] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[251:246] * PIXEL_SIZE && v_count < i_worm_y[251:246] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (42 < i_size && h_count >= i_worm_x[257:252] * PIXEL_SIZE && h_count < i_worm_x[257:252] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[257:252] * PIXEL_SIZE && v_count < i_worm_y[257:252] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (43 < i_size && h_count >= i_worm_x[263:258] * PIXEL_SIZE && h_count < i_worm_x[263:258] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[263:258] * PIXEL_SIZE && v_count < i_worm_y[263:258] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (44 < i_size && h_count >= i_worm_x[269:264] * PIXEL_SIZE && h_count < i_worm_x[269:264] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[269:264] * PIXEL_SIZE && v_count < i_worm_y[269:264] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (45 < i_size && h_count >= i_worm_x[275:270] * PIXEL_SIZE && h_count < i_worm_x[275:270] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[275:270] * PIXEL_SIZE && v_count < i_worm_y[275:270] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (46 < i_size && h_count >= i_worm_x[281:276] * PIXEL_SIZE && h_count < i_worm_x[281:276] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[281:276] * PIXEL_SIZE && v_count < i_worm_y[281:276] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (47 < i_size && h_count >= i_worm_x[287:282] * PIXEL_SIZE && h_count < i_worm_x[287:282] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[287:282] * PIXEL_SIZE && v_count < i_worm_y[287:282] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (48 < i_size && h_count >= i_worm_x[293:288] * PIXEL_SIZE && h_count < i_worm_x[293:288] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[293:288] * PIXEL_SIZE && v_count < i_worm_y[293:288] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (49 < i_size && h_count >= i_worm_x[299:294] * PIXEL_SIZE && h_count < i_worm_x[299:294] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[299:294] * PIXEL_SIZE && v_count < i_worm_y[299:294] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (50 < i_size && h_count >= i_worm_x[305:300] * PIXEL_SIZE && h_count < i_worm_x[305:300] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[305:300] * PIXEL_SIZE && v_count < i_worm_y[305:300] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (51 < i_size && h_count >= i_worm_x[311:306] * PIXEL_SIZE && h_count < i_worm_x[311:306] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[311:306] * PIXEL_SIZE && v_count < i_worm_y[311:306] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (52 < i_size && h_count >= i_worm_x[317:312] * PIXEL_SIZE && h_count < i_worm_x[317:312] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[317:312] * PIXEL_SIZE && v_count < i_worm_y[317:312] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (53 < i_size && h_count >= i_worm_x[323:318] * PIXEL_SIZE && h_count < i_worm_x[323:318] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[323:318] * PIXEL_SIZE && v_count < i_worm_y[323:318] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (54 < i_size && h_count >= i_worm_x[329:324] * PIXEL_SIZE && h_count < i_worm_x[329:324] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[329:324] * PIXEL_SIZE && v_count < i_worm_y[329:324] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (55 < i_size && h_count >= i_worm_x[335:330] * PIXEL_SIZE && h_count < i_worm_x[335:330] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[335:330] * PIXEL_SIZE && v_count < i_worm_y[335:330] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (56 < i_size && h_count >= i_worm_x[341:336] * PIXEL_SIZE && h_count < i_worm_x[341:336] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[341:336] * PIXEL_SIZE && v_count < i_worm_y[341:336] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (57 < i_size && h_count >= i_worm_x[347:342] * PIXEL_SIZE && h_count < i_worm_x[347:342] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[347:342] * PIXEL_SIZE && v_count < i_worm_y[347:342] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (58 < i_size && h_count >= i_worm_x[353:348] * PIXEL_SIZE && h_count < i_worm_x[353:348] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[353:348] * PIXEL_SIZE && v_count < i_worm_y[353:348] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (59 < i_size && h_count >= i_worm_x[359:354] * PIXEL_SIZE && h_count < i_worm_x[359:354] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[359:354] * PIXEL_SIZE && v_count < i_worm_y[359:354] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (60 < i_size && h_count >= i_worm_x[365:360] * PIXEL_SIZE && h_count < i_worm_x[365:360] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[365:360] * PIXEL_SIZE && v_count < i_worm_y[365:360] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (61 < i_size && h_count >= i_worm_x[371:366] * PIXEL_SIZE && h_count < i_worm_x[371:366] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[371:366] * PIXEL_SIZE && v_count < i_worm_y[371:366] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (62 < i_size && h_count >= i_worm_x[377:372] * PIXEL_SIZE && h_count < i_worm_x[377:372] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[377:372] * PIXEL_SIZE && v_count < i_worm_y[377:372] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (63 < i_size && h_count >= i_worm_x[383:378] * PIXEL_SIZE && h_count < i_worm_x[383:378] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[383:378] * PIXEL_SIZE && v_count < i_worm_y[383:378] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (64 < i_size && h_count >= i_worm_x[389:384] * PIXEL_SIZE && h_count < i_worm_x[389:384] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[389:384] * PIXEL_SIZE && v_count < i_worm_y[389:384] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (65 < i_size && h_count >= i_worm_x[395:390] * PIXEL_SIZE && h_count < i_worm_x[395:390] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[395:390] * PIXEL_SIZE && v_count < i_worm_y[395:390] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (66 < i_size && h_count >= i_worm_x[401:396] * PIXEL_SIZE && h_count < i_worm_x[401:396] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[401:396] * PIXEL_SIZE && v_count < i_worm_y[401:396] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (67 < i_size && h_count >= i_worm_x[407:402] * PIXEL_SIZE && h_count < i_worm_x[407:402] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[407:402] * PIXEL_SIZE && v_count < i_worm_y[407:402] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (68 < i_size && h_count >= i_worm_x[413:408] * PIXEL_SIZE && h_count < i_worm_x[413:408] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[413:408] * PIXEL_SIZE && v_count < i_worm_y[413:408] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (69 < i_size && h_count >= i_worm_x[419:414] * PIXEL_SIZE && h_count < i_worm_x[419:414] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[419:414] * PIXEL_SIZE && v_count < i_worm_y[419:414] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (70 < i_size && h_count >= i_worm_x[425:420] * PIXEL_SIZE && h_count < i_worm_x[425:420] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[425:420] * PIXEL_SIZE && v_count < i_worm_y[425:420] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (71 < i_size && h_count >= i_worm_x[431:426] * PIXEL_SIZE && h_count < i_worm_x[431:426] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[431:426] * PIXEL_SIZE && v_count < i_worm_y[431:426] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (72 < i_size && h_count >= i_worm_x[437:432] * PIXEL_SIZE && h_count < i_worm_x[437:432] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[437:432] * PIXEL_SIZE && v_count < i_worm_y[437:432] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (73 < i_size && h_count >= i_worm_x[443:438] * PIXEL_SIZE && h_count < i_worm_x[443:438] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[443:438] * PIXEL_SIZE && v_count < i_worm_y[443:438] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (74 < i_size && h_count >= i_worm_x[449:444] * PIXEL_SIZE && h_count < i_worm_x[449:444] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[449:444] * PIXEL_SIZE && v_count < i_worm_y[449:444] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (75 < i_size && h_count >= i_worm_x[455:450] * PIXEL_SIZE && h_count < i_worm_x[455:450] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[455:450] * PIXEL_SIZE && v_count < i_worm_y[455:450] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (76 < i_size && h_count >= i_worm_x[461:456] * PIXEL_SIZE && h_count < i_worm_x[461:456] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[461:456] * PIXEL_SIZE && v_count < i_worm_y[461:456] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (77 < i_size && h_count >= i_worm_x[467:462] * PIXEL_SIZE && h_count < i_worm_x[467:462] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[467:462] * PIXEL_SIZE && v_count < i_worm_y[467:462] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (78 < i_size && h_count >= i_worm_x[473:468] * PIXEL_SIZE && h_count < i_worm_x[473:468] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[473:468] * PIXEL_SIZE && v_count < i_worm_y[473:468] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (79 < i_size && h_count >= i_worm_x[479:474] * PIXEL_SIZE && h_count < i_worm_x[479:474] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[479:474] * PIXEL_SIZE && v_count < i_worm_y[479:474] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (80 < i_size && h_count >= i_worm_x[485:480] * PIXEL_SIZE && h_count < i_worm_x[485:480] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[485:480] * PIXEL_SIZE && v_count < i_worm_y[485:480] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (81 < i_size && h_count >= i_worm_x[491:486] * PIXEL_SIZE && h_count < i_worm_x[491:486] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[491:486] * PIXEL_SIZE && v_count < i_worm_y[491:486] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (82 < i_size && h_count >= i_worm_x[497:492] * PIXEL_SIZE && h_count < i_worm_x[497:492] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[497:492] * PIXEL_SIZE && v_count < i_worm_y[497:492] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (83 < i_size && h_count >= i_worm_x[503:498] * PIXEL_SIZE && h_count < i_worm_x[503:498] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[503:498] * PIXEL_SIZE && v_count < i_worm_y[503:498] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (84 < i_size && h_count >= i_worm_x[509:504] * PIXEL_SIZE && h_count < i_worm_x[509:504] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[509:504] * PIXEL_SIZE && v_count < i_worm_y[509:504] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (85 < i_size && h_count >= i_worm_x[515:510] * PIXEL_SIZE && h_count < i_worm_x[515:510] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[515:510] * PIXEL_SIZE && v_count < i_worm_y[515:510] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (86 < i_size && h_count >= i_worm_x[521:516] * PIXEL_SIZE && h_count < i_worm_x[521:516] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[521:516] * PIXEL_SIZE && v_count < i_worm_y[521:516] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (87 < i_size && h_count >= i_worm_x[527:522] * PIXEL_SIZE && h_count < i_worm_x[527:522] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[527:522] * PIXEL_SIZE && v_count < i_worm_y[527:522] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (88 < i_size && h_count >= i_worm_x[533:528] * PIXEL_SIZE && h_count < i_worm_x[533:528] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[533:528] * PIXEL_SIZE && v_count < i_worm_y[533:528] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (89 < i_size && h_count >= i_worm_x[539:534] * PIXEL_SIZE && h_count < i_worm_x[539:534] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[539:534] * PIXEL_SIZE && v_count < i_worm_y[539:534] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (90 < i_size && h_count >= i_worm_x[545:540] * PIXEL_SIZE && h_count < i_worm_x[545:540] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[545:540] * PIXEL_SIZE && v_count < i_worm_y[545:540] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (91 < i_size && h_count >= i_worm_x[551:546] * PIXEL_SIZE && h_count < i_worm_x[551:546] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[551:546] * PIXEL_SIZE && v_count < i_worm_y[551:546] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (92 < i_size && h_count >= i_worm_x[557:552] * PIXEL_SIZE && h_count < i_worm_x[557:552] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[557:552] * PIXEL_SIZE && v_count < i_worm_y[557:552] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (93 < i_size && h_count >= i_worm_x[563:558] * PIXEL_SIZE && h_count < i_worm_x[563:558] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[563:558] * PIXEL_SIZE && v_count < i_worm_y[563:558] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (94 < i_size && h_count >= i_worm_x[569:564] * PIXEL_SIZE && h_count < i_worm_x[569:564] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[569:564] * PIXEL_SIZE && v_count < i_worm_y[569:564] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (95 < i_size && h_count >= i_worm_x[575:570] * PIXEL_SIZE && h_count < i_worm_x[575:570] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[575:570] * PIXEL_SIZE && v_count < i_worm_y[575:570] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (96 < i_size && h_count >= i_worm_x[581:576] * PIXEL_SIZE && h_count < i_worm_x[581:576] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[581:576] * PIXEL_SIZE && v_count < i_worm_y[581:576] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (97 < i_size && h_count >= i_worm_x[587:582] * PIXEL_SIZE && h_count < i_worm_x[587:582] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[587:582] * PIXEL_SIZE && v_count < i_worm_y[587:582] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (98 < i_size && h_count >= i_worm_x[593:588] * PIXEL_SIZE && h_count < i_worm_x[593:588] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[593:588] * PIXEL_SIZE && v_count < i_worm_y[593:588] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (99 < i_size && h_count >= i_worm_x[599:594] * PIXEL_SIZE && h_count < i_worm_x[599:594] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[599:594] * PIXEL_SIZE && v_count < i_worm_y[599:594] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (100 < i_size && h_count >= i_worm_x[605:600] * PIXEL_SIZE && h_count < i_worm_x[605:600] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[605:600] * PIXEL_SIZE && v_count < i_worm_y[605:600] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (101 < i_size && h_count >= i_worm_x[611:606] * PIXEL_SIZE && h_count < i_worm_x[611:606] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[611:606] * PIXEL_SIZE && v_count < i_worm_y[611:606] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (102 < i_size && h_count >= i_worm_x[617:612] * PIXEL_SIZE && h_count < i_worm_x[617:612] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[617:612] * PIXEL_SIZE && v_count < i_worm_y[617:612] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (103 < i_size && h_count >= i_worm_x[623:618] * PIXEL_SIZE && h_count < i_worm_x[623:618] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[623:618] * PIXEL_SIZE && v_count < i_worm_y[623:618] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (104 < i_size && h_count >= i_worm_x[629:624] * PIXEL_SIZE && h_count < i_worm_x[629:624] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[629:624] * PIXEL_SIZE && v_count < i_worm_y[629:624] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (105 < i_size && h_count >= i_worm_x[635:630] * PIXEL_SIZE && h_count < i_worm_x[635:630] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[635:630] * PIXEL_SIZE && v_count < i_worm_y[635:630] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (106 < i_size && h_count >= i_worm_x[641:636] * PIXEL_SIZE && h_count < i_worm_x[641:636] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[641:636] * PIXEL_SIZE && v_count < i_worm_y[641:636] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (107 < i_size && h_count >= i_worm_x[647:642] * PIXEL_SIZE && h_count < i_worm_x[647:642] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[647:642] * PIXEL_SIZE && v_count < i_worm_y[647:642] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (108 < i_size && h_count >= i_worm_x[653:648] * PIXEL_SIZE && h_count < i_worm_x[653:648] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[653:648] * PIXEL_SIZE && v_count < i_worm_y[653:648] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (109 < i_size && h_count >= i_worm_x[659:654] * PIXEL_SIZE && h_count < i_worm_x[659:654] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[659:654] * PIXEL_SIZE && v_count < i_worm_y[659:654] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (110 < i_size && h_count >= i_worm_x[665:660] * PIXEL_SIZE && h_count < i_worm_x[665:660] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[665:660] * PIXEL_SIZE && v_count < i_worm_y[665:660] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (111 < i_size && h_count >= i_worm_x[671:666] * PIXEL_SIZE && h_count < i_worm_x[671:666] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[671:666] * PIXEL_SIZE && v_count < i_worm_y[671:666] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (112 < i_size && h_count >= i_worm_x[677:672] * PIXEL_SIZE && h_count < i_worm_x[677:672] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[677:672] * PIXEL_SIZE && v_count < i_worm_y[677:672] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (113 < i_size && h_count >= i_worm_x[683:678] * PIXEL_SIZE && h_count < i_worm_x[683:678] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[683:678] * PIXEL_SIZE && v_count < i_worm_y[683:678] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (114 < i_size && h_count >= i_worm_x[689:684] * PIXEL_SIZE && h_count < i_worm_x[689:684] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[689:684] * PIXEL_SIZE && v_count < i_worm_y[689:684] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (115 < i_size && h_count >= i_worm_x[695:690] * PIXEL_SIZE && h_count < i_worm_x[695:690] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[695:690] * PIXEL_SIZE && v_count < i_worm_y[695:690] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (116 < i_size && h_count >= i_worm_x[701:696] * PIXEL_SIZE && h_count < i_worm_x[701:696] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[701:696] * PIXEL_SIZE && v_count < i_worm_y[701:696] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (117 < i_size && h_count >= i_worm_x[707:702] * PIXEL_SIZE && h_count < i_worm_x[707:702] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[707:702] * PIXEL_SIZE && v_count < i_worm_y[707:702] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (118 < i_size && h_count >= i_worm_x[713:708] * PIXEL_SIZE && h_count < i_worm_x[713:708] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[713:708] * PIXEL_SIZE && v_count < i_worm_y[713:708] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (119 < i_size && h_count >= i_worm_x[719:714] * PIXEL_SIZE && h_count < i_worm_x[719:714] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[719:714] * PIXEL_SIZE && v_count < i_worm_y[719:714] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (120 < i_size && h_count >= i_worm_x[725:720] * PIXEL_SIZE && h_count < i_worm_x[725:720] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[725:720] * PIXEL_SIZE && v_count < i_worm_y[725:720] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (121 < i_size && h_count >= i_worm_x[731:726] * PIXEL_SIZE && h_count < i_worm_x[731:726] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[731:726] * PIXEL_SIZE && v_count < i_worm_y[731:726] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (122 < i_size && h_count >= i_worm_x[737:732] * PIXEL_SIZE && h_count < i_worm_x[737:732] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[737:732] * PIXEL_SIZE && v_count < i_worm_y[737:732] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (123 < i_size && h_count >= i_worm_x[743:738] * PIXEL_SIZE && h_count < i_worm_x[743:738] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[743:738] * PIXEL_SIZE && v_count < i_worm_y[743:738] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (124 < i_size && h_count >= i_worm_x[749:744] * PIXEL_SIZE && h_count < i_worm_x[749:744] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[749:744] * PIXEL_SIZE && v_count < i_worm_y[749:744] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (125 < i_size && h_count >= i_worm_x[755:750] * PIXEL_SIZE && h_count < i_worm_x[755:750] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[755:750] * PIXEL_SIZE && v_count < i_worm_y[755:750] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (126 < i_size && h_count >= i_worm_x[761:756] * PIXEL_SIZE && h_count < i_worm_x[761:756] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[761:756] * PIXEL_SIZE && v_count < i_worm_y[761:756] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (127 < i_size && h_count >= i_worm_x[767:762] * PIXEL_SIZE && h_count < i_worm_x[767:762] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[767:762] * PIXEL_SIZE && v_count < i_worm_y[767:762] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (128 < i_size && h_count >= i_worm_x[773:768] * PIXEL_SIZE && h_count < i_worm_x[773:768] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[773:768] * PIXEL_SIZE && v_count < i_worm_y[773:768] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (129 < i_size && h_count >= i_worm_x[779:774] * PIXEL_SIZE && h_count < i_worm_x[779:774] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[779:774] * PIXEL_SIZE && v_count < i_worm_y[779:774] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (130 < i_size && h_count >= i_worm_x[785:780] * PIXEL_SIZE && h_count < i_worm_x[785:780] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[785:780] * PIXEL_SIZE && v_count < i_worm_y[785:780] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (131 < i_size && h_count >= i_worm_x[791:786] * PIXEL_SIZE && h_count < i_worm_x[791:786] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[791:786] * PIXEL_SIZE && v_count < i_worm_y[791:786] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (132 < i_size && h_count >= i_worm_x[797:792] * PIXEL_SIZE && h_count < i_worm_x[797:792] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[797:792] * PIXEL_SIZE && v_count < i_worm_y[797:792] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (133 < i_size && h_count >= i_worm_x[803:798] * PIXEL_SIZE && h_count < i_worm_x[803:798] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[803:798] * PIXEL_SIZE && v_count < i_worm_y[803:798] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (134 < i_size && h_count >= i_worm_x[809:804] * PIXEL_SIZE && h_count < i_worm_x[809:804] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[809:804] * PIXEL_SIZE && v_count < i_worm_y[809:804] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (135 < i_size && h_count >= i_worm_x[815:810] * PIXEL_SIZE && h_count < i_worm_x[815:810] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[815:810] * PIXEL_SIZE && v_count < i_worm_y[815:810] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (136 < i_size && h_count >= i_worm_x[821:816] * PIXEL_SIZE && h_count < i_worm_x[821:816] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[821:816] * PIXEL_SIZE && v_count < i_worm_y[821:816] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (137 < i_size && h_count >= i_worm_x[827:822] * PIXEL_SIZE && h_count < i_worm_x[827:822] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[827:822] * PIXEL_SIZE && v_count < i_worm_y[827:822] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (138 < i_size && h_count >= i_worm_x[833:828] * PIXEL_SIZE && h_count < i_worm_x[833:828] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[833:828] * PIXEL_SIZE && v_count < i_worm_y[833:828] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (139 < i_size && h_count >= i_worm_x[839:834] * PIXEL_SIZE && h_count < i_worm_x[839:834] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[839:834] * PIXEL_SIZE && v_count < i_worm_y[839:834] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (140 < i_size && h_count >= i_worm_x[845:840] * PIXEL_SIZE && h_count < i_worm_x[845:840] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[845:840] * PIXEL_SIZE && v_count < i_worm_y[845:840] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (141 < i_size && h_count >= i_worm_x[851:846] * PIXEL_SIZE && h_count < i_worm_x[851:846] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[851:846] * PIXEL_SIZE && v_count < i_worm_y[851:846] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (142 < i_size && h_count >= i_worm_x[857:852] * PIXEL_SIZE && h_count < i_worm_x[857:852] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[857:852] * PIXEL_SIZE && v_count < i_worm_y[857:852] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (143 < i_size && h_count >= i_worm_x[863:858] * PIXEL_SIZE && h_count < i_worm_x[863:858] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[863:858] * PIXEL_SIZE && v_count < i_worm_y[863:858] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (144 < i_size && h_count >= i_worm_x[869:864] * PIXEL_SIZE && h_count < i_worm_x[869:864] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[869:864] * PIXEL_SIZE && v_count < i_worm_y[869:864] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (145 < i_size && h_count >= i_worm_x[875:870] * PIXEL_SIZE && h_count < i_worm_x[875:870] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[875:870] * PIXEL_SIZE && v_count < i_worm_y[875:870] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (146 < i_size && h_count >= i_worm_x[881:876] * PIXEL_SIZE && h_count < i_worm_x[881:876] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[881:876] * PIXEL_SIZE && v_count < i_worm_y[881:876] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (147 < i_size && h_count >= i_worm_x[887:882] * PIXEL_SIZE && h_count < i_worm_x[887:882] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[887:882] * PIXEL_SIZE && v_count < i_worm_y[887:882] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (148 < i_size && h_count >= i_worm_x[893:888] * PIXEL_SIZE && h_count < i_worm_x[893:888] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[893:888] * PIXEL_SIZE && v_count < i_worm_y[893:888] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (149 < i_size && h_count >= i_worm_x[899:894] * PIXEL_SIZE && h_count < i_worm_x[899:894] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[899:894] * PIXEL_SIZE && v_count < i_worm_y[899:894] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (150 < i_size && h_count >= i_worm_x[905:900] * PIXEL_SIZE && h_count < i_worm_x[905:900] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[905:900] * PIXEL_SIZE && v_count < i_worm_y[905:900] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (151 < i_size && h_count >= i_worm_x[911:906] * PIXEL_SIZE && h_count < i_worm_x[911:906] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[911:906] * PIXEL_SIZE && v_count < i_worm_y[911:906] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (152 < i_size && h_count >= i_worm_x[917:912] * PIXEL_SIZE && h_count < i_worm_x[917:912] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[917:912] * PIXEL_SIZE && v_count < i_worm_y[917:912] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (153 < i_size && h_count >= i_worm_x[923:918] * PIXEL_SIZE && h_count < i_worm_x[923:918] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[923:918] * PIXEL_SIZE && v_count < i_worm_y[923:918] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (154 < i_size && h_count >= i_worm_x[929:924] * PIXEL_SIZE && h_count < i_worm_x[929:924] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[929:924] * PIXEL_SIZE && v_count < i_worm_y[929:924] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (155 < i_size && h_count >= i_worm_x[935:930] * PIXEL_SIZE && h_count < i_worm_x[935:930] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[935:930] * PIXEL_SIZE && v_count < i_worm_y[935:930] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (156 < i_size && h_count >= i_worm_x[941:936] * PIXEL_SIZE && h_count < i_worm_x[941:936] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[941:936] * PIXEL_SIZE && v_count < i_worm_y[941:936] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (157 < i_size && h_count >= i_worm_x[947:942] * PIXEL_SIZE && h_count < i_worm_x[947:942] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[947:942] * PIXEL_SIZE && v_count < i_worm_y[947:942] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (158 < i_size && h_count >= i_worm_x[953:948] * PIXEL_SIZE && h_count < i_worm_x[953:948] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[953:948] * PIXEL_SIZE && v_count < i_worm_y[953:948] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (159 < i_size && h_count >= i_worm_x[959:954] * PIXEL_SIZE && h_count < i_worm_x[959:954] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[959:954] * PIXEL_SIZE && v_count < i_worm_y[959:954] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (160 < i_size && h_count >= i_worm_x[965:960] * PIXEL_SIZE && h_count < i_worm_x[965:960] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[965:960] * PIXEL_SIZE && v_count < i_worm_y[965:960] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (161 < i_size && h_count >= i_worm_x[971:966] * PIXEL_SIZE && h_count < i_worm_x[971:966] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[971:966] * PIXEL_SIZE && v_count < i_worm_y[971:966] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (162 < i_size && h_count >= i_worm_x[977:972] * PIXEL_SIZE && h_count < i_worm_x[977:972] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[977:972] * PIXEL_SIZE && v_count < i_worm_y[977:972] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (163 < i_size && h_count >= i_worm_x[983:978] * PIXEL_SIZE && h_count < i_worm_x[983:978] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[983:978] * PIXEL_SIZE && v_count < i_worm_y[983:978] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (164 < i_size && h_count >= i_worm_x[989:984] * PIXEL_SIZE && h_count < i_worm_x[989:984] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[989:984] * PIXEL_SIZE && v_count < i_worm_y[989:984] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (165 < i_size && h_count >= i_worm_x[995:990] * PIXEL_SIZE && h_count < i_worm_x[995:990] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[995:990] * PIXEL_SIZE && v_count < i_worm_y[995:990] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (166 < i_size && h_count >= i_worm_x[1001:996] * PIXEL_SIZE && h_count < i_worm_x[1001:996] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1001:996] * PIXEL_SIZE && v_count < i_worm_y[1001:996] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (167 < i_size && h_count >= i_worm_x[1007:1002] * PIXEL_SIZE && h_count < i_worm_x[1007:1002] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1007:1002] * PIXEL_SIZE && v_count < i_worm_y[1007:1002] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (168 < i_size && h_count >= i_worm_x[1013:1008] * PIXEL_SIZE && h_count < i_worm_x[1013:1008] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1013:1008] * PIXEL_SIZE && v_count < i_worm_y[1013:1008] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (169 < i_size && h_count >= i_worm_x[1019:1014] * PIXEL_SIZE && h_count < i_worm_x[1019:1014] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1019:1014] * PIXEL_SIZE && v_count < i_worm_y[1019:1014] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (170 < i_size && h_count >= i_worm_x[1025:1020] * PIXEL_SIZE && h_count < i_worm_x[1025:1020] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1025:1020] * PIXEL_SIZE && v_count < i_worm_y[1025:1020] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (171 < i_size && h_count >= i_worm_x[1031:1026] * PIXEL_SIZE && h_count < i_worm_x[1031:1026] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1031:1026] * PIXEL_SIZE && v_count < i_worm_y[1031:1026] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (172 < i_size && h_count >= i_worm_x[1037:1032] * PIXEL_SIZE && h_count < i_worm_x[1037:1032] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1037:1032] * PIXEL_SIZE && v_count < i_worm_y[1037:1032] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (173 < i_size && h_count >= i_worm_x[1043:1038] * PIXEL_SIZE && h_count < i_worm_x[1043:1038] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1043:1038] * PIXEL_SIZE && v_count < i_worm_y[1043:1038] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (174 < i_size && h_count >= i_worm_x[1049:1044] * PIXEL_SIZE && h_count < i_worm_x[1049:1044] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1049:1044] * PIXEL_SIZE && v_count < i_worm_y[1049:1044] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (175 < i_size && h_count >= i_worm_x[1055:1050] * PIXEL_SIZE && h_count < i_worm_x[1055:1050] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1055:1050] * PIXEL_SIZE && v_count < i_worm_y[1055:1050] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (176 < i_size && h_count >= i_worm_x[1061:1056] * PIXEL_SIZE && h_count < i_worm_x[1061:1056] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1061:1056] * PIXEL_SIZE && v_count < i_worm_y[1061:1056] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (177 < i_size && h_count >= i_worm_x[1067:1062] * PIXEL_SIZE && h_count < i_worm_x[1067:1062] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1067:1062] * PIXEL_SIZE && v_count < i_worm_y[1067:1062] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (178 < i_size && h_count >= i_worm_x[1073:1068] * PIXEL_SIZE && h_count < i_worm_x[1073:1068] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1073:1068] * PIXEL_SIZE && v_count < i_worm_y[1073:1068] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (179 < i_size && h_count >= i_worm_x[1079:1074] * PIXEL_SIZE && h_count < i_worm_x[1079:1074] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1079:1074] * PIXEL_SIZE && v_count < i_worm_y[1079:1074] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (180 < i_size && h_count >= i_worm_x[1085:1080] * PIXEL_SIZE && h_count < i_worm_x[1085:1080] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1085:1080] * PIXEL_SIZE && v_count < i_worm_y[1085:1080] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (181 < i_size && h_count >= i_worm_x[1091:1086] * PIXEL_SIZE && h_count < i_worm_x[1091:1086] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1091:1086] * PIXEL_SIZE && v_count < i_worm_y[1091:1086] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (182 < i_size && h_count >= i_worm_x[1097:1092] * PIXEL_SIZE && h_count < i_worm_x[1097:1092] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1097:1092] * PIXEL_SIZE && v_count < i_worm_y[1097:1092] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (183 < i_size && h_count >= i_worm_x[1103:1098] * PIXEL_SIZE && h_count < i_worm_x[1103:1098] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1103:1098] * PIXEL_SIZE && v_count < i_worm_y[1103:1098] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (184 < i_size && h_count >= i_worm_x[1109:1104] * PIXEL_SIZE && h_count < i_worm_x[1109:1104] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1109:1104] * PIXEL_SIZE && v_count < i_worm_y[1109:1104] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (185 < i_size && h_count >= i_worm_x[1115:1110] * PIXEL_SIZE && h_count < i_worm_x[1115:1110] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1115:1110] * PIXEL_SIZE && v_count < i_worm_y[1115:1110] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (186 < i_size && h_count >= i_worm_x[1121:1116] * PIXEL_SIZE && h_count < i_worm_x[1121:1116] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1121:1116] * PIXEL_SIZE && v_count < i_worm_y[1121:1116] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (187 < i_size && h_count >= i_worm_x[1127:1122] * PIXEL_SIZE && h_count < i_worm_x[1127:1122] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1127:1122] * PIXEL_SIZE && v_count < i_worm_y[1127:1122] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (188 < i_size && h_count >= i_worm_x[1133:1128] * PIXEL_SIZE && h_count < i_worm_x[1133:1128] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1133:1128] * PIXEL_SIZE && v_count < i_worm_y[1133:1128] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (189 < i_size && h_count >= i_worm_x[1139:1134] * PIXEL_SIZE && h_count < i_worm_x[1139:1134] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1139:1134] * PIXEL_SIZE && v_count < i_worm_y[1139:1134] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (190 < i_size && h_count >= i_worm_x[1145:1140] * PIXEL_SIZE && h_count < i_worm_x[1145:1140] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1145:1140] * PIXEL_SIZE && v_count < i_worm_y[1145:1140] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (191 < i_size && h_count >= i_worm_x[1151:1146] * PIXEL_SIZE && h_count < i_worm_x[1151:1146] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1151:1146] * PIXEL_SIZE && v_count < i_worm_y[1151:1146] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (192 < i_size && h_count >= i_worm_x[1157:1152] * PIXEL_SIZE && h_count < i_worm_x[1157:1152] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1157:1152] * PIXEL_SIZE && v_count < i_worm_y[1157:1152] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (193 < i_size && h_count >= i_worm_x[1163:1158] * PIXEL_SIZE && h_count < i_worm_x[1163:1158] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1163:1158] * PIXEL_SIZE && v_count < i_worm_y[1163:1158] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (194 < i_size && h_count >= i_worm_x[1169:1164] * PIXEL_SIZE && h_count < i_worm_x[1169:1164] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1169:1164] * PIXEL_SIZE && v_count < i_worm_y[1169:1164] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (195 < i_size && h_count >= i_worm_x[1175:1170] * PIXEL_SIZE && h_count < i_worm_x[1175:1170] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1175:1170] * PIXEL_SIZE && v_count < i_worm_y[1175:1170] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (196 < i_size && h_count >= i_worm_x[1181:1176] * PIXEL_SIZE && h_count < i_worm_x[1181:1176] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1181:1176] * PIXEL_SIZE && v_count < i_worm_y[1181:1176] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (197 < i_size && h_count >= i_worm_x[1187:1182] * PIXEL_SIZE && h_count < i_worm_x[1187:1182] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1187:1182] * PIXEL_SIZE && v_count < i_worm_y[1187:1182] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (198 < i_size && h_count >= i_worm_x[1193:1188] * PIXEL_SIZE && h_count < i_worm_x[1193:1188] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1193:1188] * PIXEL_SIZE && v_count < i_worm_y[1193:1188] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (199 < i_size && h_count >= i_worm_x[1199:1194] * PIXEL_SIZE && h_count < i_worm_x[1199:1194] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1199:1194] * PIXEL_SIZE && v_count < i_worm_y[1199:1194] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (200 < i_size && h_count >= i_worm_x[1205:1200] * PIXEL_SIZE && h_count < i_worm_x[1205:1200] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1205:1200] * PIXEL_SIZE && v_count < i_worm_y[1205:1200] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (201 < i_size && h_count >= i_worm_x[1211:1206] * PIXEL_SIZE && h_count < i_worm_x[1211:1206] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1211:1206] * PIXEL_SIZE && v_count < i_worm_y[1211:1206] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (202 < i_size && h_count >= i_worm_x[1217:1212] * PIXEL_SIZE && h_count < i_worm_x[1217:1212] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1217:1212] * PIXEL_SIZE && v_count < i_worm_y[1217:1212] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (203 < i_size && h_count >= i_worm_x[1223:1218] * PIXEL_SIZE && h_count < i_worm_x[1223:1218] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1223:1218] * PIXEL_SIZE && v_count < i_worm_y[1223:1218] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (204 < i_size && h_count >= i_worm_x[1229:1224] * PIXEL_SIZE && h_count < i_worm_x[1229:1224] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1229:1224] * PIXEL_SIZE && v_count < i_worm_y[1229:1224] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (205 < i_size && h_count >= i_worm_x[1235:1230] * PIXEL_SIZE && h_count < i_worm_x[1235:1230] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1235:1230] * PIXEL_SIZE && v_count < i_worm_y[1235:1230] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (206 < i_size && h_count >= i_worm_x[1241:1236] * PIXEL_SIZE && h_count < i_worm_x[1241:1236] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1241:1236] * PIXEL_SIZE && v_count < i_worm_y[1241:1236] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (207 < i_size && h_count >= i_worm_x[1247:1242] * PIXEL_SIZE && h_count < i_worm_x[1247:1242] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1247:1242] * PIXEL_SIZE && v_count < i_worm_y[1247:1242] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (208 < i_size && h_count >= i_worm_x[1253:1248] * PIXEL_SIZE && h_count < i_worm_x[1253:1248] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1253:1248] * PIXEL_SIZE && v_count < i_worm_y[1253:1248] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (209 < i_size && h_count >= i_worm_x[1259:1254] * PIXEL_SIZE && h_count < i_worm_x[1259:1254] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1259:1254] * PIXEL_SIZE && v_count < i_worm_y[1259:1254] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (210 < i_size && h_count >= i_worm_x[1265:1260] * PIXEL_SIZE && h_count < i_worm_x[1265:1260] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1265:1260] * PIXEL_SIZE && v_count < i_worm_y[1265:1260] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (211 < i_size && h_count >= i_worm_x[1271:1266] * PIXEL_SIZE && h_count < i_worm_x[1271:1266] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1271:1266] * PIXEL_SIZE && v_count < i_worm_y[1271:1266] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (212 < i_size && h_count >= i_worm_x[1277:1272] * PIXEL_SIZE && h_count < i_worm_x[1277:1272] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1277:1272] * PIXEL_SIZE && v_count < i_worm_y[1277:1272] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (213 < i_size && h_count >= i_worm_x[1283:1278] * PIXEL_SIZE && h_count < i_worm_x[1283:1278] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1283:1278] * PIXEL_SIZE && v_count < i_worm_y[1283:1278] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (214 < i_size && h_count >= i_worm_x[1289:1284] * PIXEL_SIZE && h_count < i_worm_x[1289:1284] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1289:1284] * PIXEL_SIZE && v_count < i_worm_y[1289:1284] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (215 < i_size && h_count >= i_worm_x[1295:1290] * PIXEL_SIZE && h_count < i_worm_x[1295:1290] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1295:1290] * PIXEL_SIZE && v_count < i_worm_y[1295:1290] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (216 < i_size && h_count >= i_worm_x[1301:1296] * PIXEL_SIZE && h_count < i_worm_x[1301:1296] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1301:1296] * PIXEL_SIZE && v_count < i_worm_y[1301:1296] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (217 < i_size && h_count >= i_worm_x[1307:1302] * PIXEL_SIZE && h_count < i_worm_x[1307:1302] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1307:1302] * PIXEL_SIZE && v_count < i_worm_y[1307:1302] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (218 < i_size && h_count >= i_worm_x[1313:1308] * PIXEL_SIZE && h_count < i_worm_x[1313:1308] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1313:1308] * PIXEL_SIZE && v_count < i_worm_y[1313:1308] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (219 < i_size && h_count >= i_worm_x[1319:1314] * PIXEL_SIZE && h_count < i_worm_x[1319:1314] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1319:1314] * PIXEL_SIZE && v_count < i_worm_y[1319:1314] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (220 < i_size && h_count >= i_worm_x[1325:1320] * PIXEL_SIZE && h_count < i_worm_x[1325:1320] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1325:1320] * PIXEL_SIZE && v_count < i_worm_y[1325:1320] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (221 < i_size && h_count >= i_worm_x[1331:1326] * PIXEL_SIZE && h_count < i_worm_x[1331:1326] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1331:1326] * PIXEL_SIZE && v_count < i_worm_y[1331:1326] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (222 < i_size && h_count >= i_worm_x[1337:1332] * PIXEL_SIZE && h_count < i_worm_x[1337:1332] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1337:1332] * PIXEL_SIZE && v_count < i_worm_y[1337:1332] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (223 < i_size && h_count >= i_worm_x[1343:1338] * PIXEL_SIZE && h_count < i_worm_x[1343:1338] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1343:1338] * PIXEL_SIZE && v_count < i_worm_y[1343:1338] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (224 < i_size && h_count >= i_worm_x[1349:1344] * PIXEL_SIZE && h_count < i_worm_x[1349:1344] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1349:1344] * PIXEL_SIZE && v_count < i_worm_y[1349:1344] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (225 < i_size && h_count >= i_worm_x[1355:1350] * PIXEL_SIZE && h_count < i_worm_x[1355:1350] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1355:1350] * PIXEL_SIZE && v_count < i_worm_y[1355:1350] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (226 < i_size && h_count >= i_worm_x[1361:1356] * PIXEL_SIZE && h_count < i_worm_x[1361:1356] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1361:1356] * PIXEL_SIZE && v_count < i_worm_y[1361:1356] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (227 < i_size && h_count >= i_worm_x[1367:1362] * PIXEL_SIZE && h_count < i_worm_x[1367:1362] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1367:1362] * PIXEL_SIZE && v_count < i_worm_y[1367:1362] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (228 < i_size && h_count >= i_worm_x[1373:1368] * PIXEL_SIZE && h_count < i_worm_x[1373:1368] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1373:1368] * PIXEL_SIZE && v_count < i_worm_y[1373:1368] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (229 < i_size && h_count >= i_worm_x[1379:1374] * PIXEL_SIZE && h_count < i_worm_x[1379:1374] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1379:1374] * PIXEL_SIZE && v_count < i_worm_y[1379:1374] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (230 < i_size && h_count >= i_worm_x[1385:1380] * PIXEL_SIZE && h_count < i_worm_x[1385:1380] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1385:1380] * PIXEL_SIZE && v_count < i_worm_y[1385:1380] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (231 < i_size && h_count >= i_worm_x[1391:1386] * PIXEL_SIZE && h_count < i_worm_x[1391:1386] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1391:1386] * PIXEL_SIZE && v_count < i_worm_y[1391:1386] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (232 < i_size && h_count >= i_worm_x[1397:1392] * PIXEL_SIZE && h_count < i_worm_x[1397:1392] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1397:1392] * PIXEL_SIZE && v_count < i_worm_y[1397:1392] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (233 < i_size && h_count >= i_worm_x[1403:1398] * PIXEL_SIZE && h_count < i_worm_x[1403:1398] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1403:1398] * PIXEL_SIZE && v_count < i_worm_y[1403:1398] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (234 < i_size && h_count >= i_worm_x[1409:1404] * PIXEL_SIZE && h_count < i_worm_x[1409:1404] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1409:1404] * PIXEL_SIZE && v_count < i_worm_y[1409:1404] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (235 < i_size && h_count >= i_worm_x[1415:1410] * PIXEL_SIZE && h_count < i_worm_x[1415:1410] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1415:1410] * PIXEL_SIZE && v_count < i_worm_y[1415:1410] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (236 < i_size && h_count >= i_worm_x[1421:1416] * PIXEL_SIZE && h_count < i_worm_x[1421:1416] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1421:1416] * PIXEL_SIZE && v_count < i_worm_y[1421:1416] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (237 < i_size && h_count >= i_worm_x[1427:1422] * PIXEL_SIZE && h_count < i_worm_x[1427:1422] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1427:1422] * PIXEL_SIZE && v_count < i_worm_y[1427:1422] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (238 < i_size && h_count >= i_worm_x[1433:1428] * PIXEL_SIZE && h_count < i_worm_x[1433:1428] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1433:1428] * PIXEL_SIZE && v_count < i_worm_y[1433:1428] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (239 < i_size && h_count >= i_worm_x[1439:1434] * PIXEL_SIZE && h_count < i_worm_x[1439:1434] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1439:1434] * PIXEL_SIZE && v_count < i_worm_y[1439:1434] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (240 < i_size && h_count >= i_worm_x[1445:1440] * PIXEL_SIZE && h_count < i_worm_x[1445:1440] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1445:1440] * PIXEL_SIZE && v_count < i_worm_y[1445:1440] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (241 < i_size && h_count >= i_worm_x[1451:1446] * PIXEL_SIZE && h_count < i_worm_x[1451:1446] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1451:1446] * PIXEL_SIZE && v_count < i_worm_y[1451:1446] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (242 < i_size && h_count >= i_worm_x[1457:1452] * PIXEL_SIZE && h_count < i_worm_x[1457:1452] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1457:1452] * PIXEL_SIZE && v_count < i_worm_y[1457:1452] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (243 < i_size && h_count >= i_worm_x[1463:1458] * PIXEL_SIZE && h_count < i_worm_x[1463:1458] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1463:1458] * PIXEL_SIZE && v_count < i_worm_y[1463:1458] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (244 < i_size && h_count >= i_worm_x[1469:1464] * PIXEL_SIZE && h_count < i_worm_x[1469:1464] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1469:1464] * PIXEL_SIZE && v_count < i_worm_y[1469:1464] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (245 < i_size && h_count >= i_worm_x[1475:1470] * PIXEL_SIZE && h_count < i_worm_x[1475:1470] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1475:1470] * PIXEL_SIZE && v_count < i_worm_y[1475:1470] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (246 < i_size && h_count >= i_worm_x[1481:1476] * PIXEL_SIZE && h_count < i_worm_x[1481:1476] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1481:1476] * PIXEL_SIZE && v_count < i_worm_y[1481:1476] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (247 < i_size && h_count >= i_worm_x[1487:1482] * PIXEL_SIZE && h_count < i_worm_x[1487:1482] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1487:1482] * PIXEL_SIZE && v_count < i_worm_y[1487:1482] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (248 < i_size && h_count >= i_worm_x[1493:1488] * PIXEL_SIZE && h_count < i_worm_x[1493:1488] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1493:1488] * PIXEL_SIZE && v_count < i_worm_y[1493:1488] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (249 < i_size && h_count >= i_worm_x[1499:1494] * PIXEL_SIZE && h_count < i_worm_x[1499:1494] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1499:1494] * PIXEL_SIZE && v_count < i_worm_y[1499:1494] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (250 < i_size && h_count >= i_worm_x[1505:1500] * PIXEL_SIZE && h_count < i_worm_x[1505:1500] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1505:1500] * PIXEL_SIZE && v_count < i_worm_y[1505:1500] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (251 < i_size && h_count >= i_worm_x[1511:1506] * PIXEL_SIZE && h_count < i_worm_x[1511:1506] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1511:1506] * PIXEL_SIZE && v_count < i_worm_y[1511:1506] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (252 < i_size && h_count >= i_worm_x[1517:1512] * PIXEL_SIZE && h_count < i_worm_x[1517:1512] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1517:1512] * PIXEL_SIZE && v_count < i_worm_y[1517:1512] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (253 < i_size && h_count >= i_worm_x[1523:1518] * PIXEL_SIZE && h_count < i_worm_x[1523:1518] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1523:1518] * PIXEL_SIZE && v_count < i_worm_y[1523:1518] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (254 < i_size && h_count >= i_worm_x[1529:1524] * PIXEL_SIZE && h_count < i_worm_x[1529:1524] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1529:1524] * PIXEL_SIZE && v_count < i_worm_y[1529:1524] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (255 < i_size && h_count >= i_worm_x[1535:1530] * PIXEL_SIZE && h_count < i_worm_x[1535:1530] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1535:1530] * PIXEL_SIZE && v_count < i_worm_y[1535:1530] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (256 < i_size && h_count >= i_worm_x[1541:1536] * PIXEL_SIZE && h_count < i_worm_x[1541:1536] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1541:1536] * PIXEL_SIZE && v_count < i_worm_y[1541:1536] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (257 < i_size && h_count >= i_worm_x[1547:1542] * PIXEL_SIZE && h_count < i_worm_x[1547:1542] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1547:1542] * PIXEL_SIZE && v_count < i_worm_y[1547:1542] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (258 < i_size && h_count >= i_worm_x[1553:1548] * PIXEL_SIZE && h_count < i_worm_x[1553:1548] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1553:1548] * PIXEL_SIZE && v_count < i_worm_y[1553:1548] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (259 < i_size && h_count >= i_worm_x[1559:1554] * PIXEL_SIZE && h_count < i_worm_x[1559:1554] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1559:1554] * PIXEL_SIZE && v_count < i_worm_y[1559:1554] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (260 < i_size && h_count >= i_worm_x[1565:1560] * PIXEL_SIZE && h_count < i_worm_x[1565:1560] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1565:1560] * PIXEL_SIZE && v_count < i_worm_y[1565:1560] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (261 < i_size && h_count >= i_worm_x[1571:1566] * PIXEL_SIZE && h_count < i_worm_x[1571:1566] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1571:1566] * PIXEL_SIZE && v_count < i_worm_y[1571:1566] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (262 < i_size && h_count >= i_worm_x[1577:1572] * PIXEL_SIZE && h_count < i_worm_x[1577:1572] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1577:1572] * PIXEL_SIZE && v_count < i_worm_y[1577:1572] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (263 < i_size && h_count >= i_worm_x[1583:1578] * PIXEL_SIZE && h_count < i_worm_x[1583:1578] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1583:1578] * PIXEL_SIZE && v_count < i_worm_y[1583:1578] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (264 < i_size && h_count >= i_worm_x[1589:1584] * PIXEL_SIZE && h_count < i_worm_x[1589:1584] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1589:1584] * PIXEL_SIZE && v_count < i_worm_y[1589:1584] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (265 < i_size && h_count >= i_worm_x[1595:1590] * PIXEL_SIZE && h_count < i_worm_x[1595:1590] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1595:1590] * PIXEL_SIZE && v_count < i_worm_y[1595:1590] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (266 < i_size && h_count >= i_worm_x[1601:1596] * PIXEL_SIZE && h_count < i_worm_x[1601:1596] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1601:1596] * PIXEL_SIZE && v_count < i_worm_y[1601:1596] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (267 < i_size && h_count >= i_worm_x[1607:1602] * PIXEL_SIZE && h_count < i_worm_x[1607:1602] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1607:1602] * PIXEL_SIZE && v_count < i_worm_y[1607:1602] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (268 < i_size && h_count >= i_worm_x[1613:1608] * PIXEL_SIZE && h_count < i_worm_x[1613:1608] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1613:1608] * PIXEL_SIZE && v_count < i_worm_y[1613:1608] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (269 < i_size && h_count >= i_worm_x[1619:1614] * PIXEL_SIZE && h_count < i_worm_x[1619:1614] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1619:1614] * PIXEL_SIZE && v_count < i_worm_y[1619:1614] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (270 < i_size && h_count >= i_worm_x[1625:1620] * PIXEL_SIZE && h_count < i_worm_x[1625:1620] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1625:1620] * PIXEL_SIZE && v_count < i_worm_y[1625:1620] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (271 < i_size && h_count >= i_worm_x[1631:1626] * PIXEL_SIZE && h_count < i_worm_x[1631:1626] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1631:1626] * PIXEL_SIZE && v_count < i_worm_y[1631:1626] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (272 < i_size && h_count >= i_worm_x[1637:1632] * PIXEL_SIZE && h_count < i_worm_x[1637:1632] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1637:1632] * PIXEL_SIZE && v_count < i_worm_y[1637:1632] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (273 < i_size && h_count >= i_worm_x[1643:1638] * PIXEL_SIZE && h_count < i_worm_x[1643:1638] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1643:1638] * PIXEL_SIZE && v_count < i_worm_y[1643:1638] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (274 < i_size && h_count >= i_worm_x[1649:1644] * PIXEL_SIZE && h_count < i_worm_x[1649:1644] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1649:1644] * PIXEL_SIZE && v_count < i_worm_y[1649:1644] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (275 < i_size && h_count >= i_worm_x[1655:1650] * PIXEL_SIZE && h_count < i_worm_x[1655:1650] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1655:1650] * PIXEL_SIZE && v_count < i_worm_y[1655:1650] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (276 < i_size && h_count >= i_worm_x[1661:1656] * PIXEL_SIZE && h_count < i_worm_x[1661:1656] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1661:1656] * PIXEL_SIZE && v_count < i_worm_y[1661:1656] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (277 < i_size && h_count >= i_worm_x[1667:1662] * PIXEL_SIZE && h_count < i_worm_x[1667:1662] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1667:1662] * PIXEL_SIZE && v_count < i_worm_y[1667:1662] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (278 < i_size && h_count >= i_worm_x[1673:1668] * PIXEL_SIZE && h_count < i_worm_x[1673:1668] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1673:1668] * PIXEL_SIZE && v_count < i_worm_y[1673:1668] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (279 < i_size && h_count >= i_worm_x[1679:1674] * PIXEL_SIZE && h_count < i_worm_x[1679:1674] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1679:1674] * PIXEL_SIZE && v_count < i_worm_y[1679:1674] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (280 < i_size && h_count >= i_worm_x[1685:1680] * PIXEL_SIZE && h_count < i_worm_x[1685:1680] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1685:1680] * PIXEL_SIZE && v_count < i_worm_y[1685:1680] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (281 < i_size && h_count >= i_worm_x[1691:1686] * PIXEL_SIZE && h_count < i_worm_x[1691:1686] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1691:1686] * PIXEL_SIZE && v_count < i_worm_y[1691:1686] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (282 < i_size && h_count >= i_worm_x[1697:1692] * PIXEL_SIZE && h_count < i_worm_x[1697:1692] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1697:1692] * PIXEL_SIZE && v_count < i_worm_y[1697:1692] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (283 < i_size && h_count >= i_worm_x[1703:1698] * PIXEL_SIZE && h_count < i_worm_x[1703:1698] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1703:1698] * PIXEL_SIZE && v_count < i_worm_y[1703:1698] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (284 < i_size && h_count >= i_worm_x[1709:1704] * PIXEL_SIZE && h_count < i_worm_x[1709:1704] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1709:1704] * PIXEL_SIZE && v_count < i_worm_y[1709:1704] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (285 < i_size && h_count >= i_worm_x[1715:1710] * PIXEL_SIZE && h_count < i_worm_x[1715:1710] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1715:1710] * PIXEL_SIZE && v_count < i_worm_y[1715:1710] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (286 < i_size && h_count >= i_worm_x[1721:1716] * PIXEL_SIZE && h_count < i_worm_x[1721:1716] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1721:1716] * PIXEL_SIZE && v_count < i_worm_y[1721:1716] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (287 < i_size && h_count >= i_worm_x[1727:1722] * PIXEL_SIZE && h_count < i_worm_x[1727:1722] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1727:1722] * PIXEL_SIZE && v_count < i_worm_y[1727:1722] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (288 < i_size && h_count >= i_worm_x[1733:1728] * PIXEL_SIZE && h_count < i_worm_x[1733:1728] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1733:1728] * PIXEL_SIZE && v_count < i_worm_y[1733:1728] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (289 < i_size && h_count >= i_worm_x[1739:1734] * PIXEL_SIZE && h_count < i_worm_x[1739:1734] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1739:1734] * PIXEL_SIZE && v_count < i_worm_y[1739:1734] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (290 < i_size && h_count >= i_worm_x[1745:1740] * PIXEL_SIZE && h_count < i_worm_x[1745:1740] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1745:1740] * PIXEL_SIZE && v_count < i_worm_y[1745:1740] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (291 < i_size && h_count >= i_worm_x[1751:1746] * PIXEL_SIZE && h_count < i_worm_x[1751:1746] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1751:1746] * PIXEL_SIZE && v_count < i_worm_y[1751:1746] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (292 < i_size && h_count >= i_worm_x[1757:1752] * PIXEL_SIZE && h_count < i_worm_x[1757:1752] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1757:1752] * PIXEL_SIZE && v_count < i_worm_y[1757:1752] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (293 < i_size && h_count >= i_worm_x[1763:1758] * PIXEL_SIZE && h_count < i_worm_x[1763:1758] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1763:1758] * PIXEL_SIZE && v_count < i_worm_y[1763:1758] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (294 < i_size && h_count >= i_worm_x[1769:1764] * PIXEL_SIZE && h_count < i_worm_x[1769:1764] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1769:1764] * PIXEL_SIZE && v_count < i_worm_y[1769:1764] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (295 < i_size && h_count >= i_worm_x[1775:1770] * PIXEL_SIZE && h_count < i_worm_x[1775:1770] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1775:1770] * PIXEL_SIZE && v_count < i_worm_y[1775:1770] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (296 < i_size && h_count >= i_worm_x[1781:1776] * PIXEL_SIZE && h_count < i_worm_x[1781:1776] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1781:1776] * PIXEL_SIZE && v_count < i_worm_y[1781:1776] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (297 < i_size && h_count >= i_worm_x[1787:1782] * PIXEL_SIZE && h_count < i_worm_x[1787:1782] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1787:1782] * PIXEL_SIZE && v_count < i_worm_y[1787:1782] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (298 < i_size && h_count >= i_worm_x[1793:1788] * PIXEL_SIZE && h_count < i_worm_x[1793:1788] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1793:1788] * PIXEL_SIZE && v_count < i_worm_y[1793:1788] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (299 < i_size && h_count >= i_worm_x[1799:1794] * PIXEL_SIZE && h_count < i_worm_x[1799:1794] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1799:1794] * PIXEL_SIZE && v_count < i_worm_y[1799:1794] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (300 < i_size && h_count >= i_worm_x[1805:1800] * PIXEL_SIZE && h_count < i_worm_x[1805:1800] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1805:1800] * PIXEL_SIZE && v_count < i_worm_y[1805:1800] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (301 < i_size && h_count >= i_worm_x[1811:1806] * PIXEL_SIZE && h_count < i_worm_x[1811:1806] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1811:1806] * PIXEL_SIZE && v_count < i_worm_y[1811:1806] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (302 < i_size && h_count >= i_worm_x[1817:1812] * PIXEL_SIZE && h_count < i_worm_x[1817:1812] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1817:1812] * PIXEL_SIZE && v_count < i_worm_y[1817:1812] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (303 < i_size && h_count >= i_worm_x[1823:1818] * PIXEL_SIZE && h_count < i_worm_x[1823:1818] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1823:1818] * PIXEL_SIZE && v_count < i_worm_y[1823:1818] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (304 < i_size && h_count >= i_worm_x[1829:1824] * PIXEL_SIZE && h_count < i_worm_x[1829:1824] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1829:1824] * PIXEL_SIZE && v_count < i_worm_y[1829:1824] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (305 < i_size && h_count >= i_worm_x[1835:1830] * PIXEL_SIZE && h_count < i_worm_x[1835:1830] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1835:1830] * PIXEL_SIZE && v_count < i_worm_y[1835:1830] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (306 < i_size && h_count >= i_worm_x[1841:1836] * PIXEL_SIZE && h_count < i_worm_x[1841:1836] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1841:1836] * PIXEL_SIZE && v_count < i_worm_y[1841:1836] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (307 < i_size && h_count >= i_worm_x[1847:1842] * PIXEL_SIZE && h_count < i_worm_x[1847:1842] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1847:1842] * PIXEL_SIZE && v_count < i_worm_y[1847:1842] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (308 < i_size && h_count >= i_worm_x[1853:1848] * PIXEL_SIZE && h_count < i_worm_x[1853:1848] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1853:1848] * PIXEL_SIZE && v_count < i_worm_y[1853:1848] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (309 < i_size && h_count >= i_worm_x[1859:1854] * PIXEL_SIZE && h_count < i_worm_x[1859:1854] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1859:1854] * PIXEL_SIZE && v_count < i_worm_y[1859:1854] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (310 < i_size && h_count >= i_worm_x[1865:1860] * PIXEL_SIZE && h_count < i_worm_x[1865:1860] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1865:1860] * PIXEL_SIZE && v_count < i_worm_y[1865:1860] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (311 < i_size && h_count >= i_worm_x[1871:1866] * PIXEL_SIZE && h_count < i_worm_x[1871:1866] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1871:1866] * PIXEL_SIZE && v_count < i_worm_y[1871:1866] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (312 < i_size && h_count >= i_worm_x[1877:1872] * PIXEL_SIZE && h_count < i_worm_x[1877:1872] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1877:1872] * PIXEL_SIZE && v_count < i_worm_y[1877:1872] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (313 < i_size && h_count >= i_worm_x[1883:1878] * PIXEL_SIZE && h_count < i_worm_x[1883:1878] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1883:1878] * PIXEL_SIZE && v_count < i_worm_y[1883:1878] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (314 < i_size && h_count >= i_worm_x[1889:1884] * PIXEL_SIZE && h_count < i_worm_x[1889:1884] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1889:1884] * PIXEL_SIZE && v_count < i_worm_y[1889:1884] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (315 < i_size && h_count >= i_worm_x[1895:1890] * PIXEL_SIZE && h_count < i_worm_x[1895:1890] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1895:1890] * PIXEL_SIZE && v_count < i_worm_y[1895:1890] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (316 < i_size && h_count >= i_worm_x[1901:1896] * PIXEL_SIZE && h_count < i_worm_x[1901:1896] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1901:1896] * PIXEL_SIZE && v_count < i_worm_y[1901:1896] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (317 < i_size && h_count >= i_worm_x[1907:1902] * PIXEL_SIZE && h_count < i_worm_x[1907:1902] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1907:1902] * PIXEL_SIZE && v_count < i_worm_y[1907:1902] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (318 < i_size && h_count >= i_worm_x[1913:1908] * PIXEL_SIZE && h_count < i_worm_x[1913:1908] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1913:1908] * PIXEL_SIZE && v_count < i_worm_y[1913:1908] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (319 < i_size && h_count >= i_worm_x[1919:1914] * PIXEL_SIZE && h_count < i_worm_x[1919:1914] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1919:1914] * PIXEL_SIZE && v_count < i_worm_y[1919:1914] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (320 < i_size && h_count >= i_worm_x[1925:1920] * PIXEL_SIZE && h_count < i_worm_x[1925:1920] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1925:1920] * PIXEL_SIZE && v_count < i_worm_y[1925:1920] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (321 < i_size && h_count >= i_worm_x[1931:1926] * PIXEL_SIZE && h_count < i_worm_x[1931:1926] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1931:1926] * PIXEL_SIZE && v_count < i_worm_y[1931:1926] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (322 < i_size && h_count >= i_worm_x[1937:1932] * PIXEL_SIZE && h_count < i_worm_x[1937:1932] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1937:1932] * PIXEL_SIZE && v_count < i_worm_y[1937:1932] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (323 < i_size && h_count >= i_worm_x[1943:1938] * PIXEL_SIZE && h_count < i_worm_x[1943:1938] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1943:1938] * PIXEL_SIZE && v_count < i_worm_y[1943:1938] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (324 < i_size && h_count >= i_worm_x[1949:1944] * PIXEL_SIZE && h_count < i_worm_x[1949:1944] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1949:1944] * PIXEL_SIZE && v_count < i_worm_y[1949:1944] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (325 < i_size && h_count >= i_worm_x[1955:1950] * PIXEL_SIZE && h_count < i_worm_x[1955:1950] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1955:1950] * PIXEL_SIZE && v_count < i_worm_y[1955:1950] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (326 < i_size && h_count >= i_worm_x[1961:1956] * PIXEL_SIZE && h_count < i_worm_x[1961:1956] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1961:1956] * PIXEL_SIZE && v_count < i_worm_y[1961:1956] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (327 < i_size && h_count >= i_worm_x[1967:1962] * PIXEL_SIZE && h_count < i_worm_x[1967:1962] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1967:1962] * PIXEL_SIZE && v_count < i_worm_y[1967:1962] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (328 < i_size && h_count >= i_worm_x[1973:1968] * PIXEL_SIZE && h_count < i_worm_x[1973:1968] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1973:1968] * PIXEL_SIZE && v_count < i_worm_y[1973:1968] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (329 < i_size && h_count >= i_worm_x[1979:1974] * PIXEL_SIZE && h_count < i_worm_x[1979:1974] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1979:1974] * PIXEL_SIZE && v_count < i_worm_y[1979:1974] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (330 < i_size && h_count >= i_worm_x[1985:1980] * PIXEL_SIZE && h_count < i_worm_x[1985:1980] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1985:1980] * PIXEL_SIZE && v_count < i_worm_y[1985:1980] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (331 < i_size && h_count >= i_worm_x[1991:1986] * PIXEL_SIZE && h_count < i_worm_x[1991:1986] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1991:1986] * PIXEL_SIZE && v_count < i_worm_y[1991:1986] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (332 < i_size && h_count >= i_worm_x[1997:1992] * PIXEL_SIZE && h_count < i_worm_x[1997:1992] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[1997:1992] * PIXEL_SIZE && v_count < i_worm_y[1997:1992] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (333 < i_size && h_count >= i_worm_x[2003:1998] * PIXEL_SIZE && h_count < i_worm_x[2003:1998] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2003:1998] * PIXEL_SIZE && v_count < i_worm_y[2003:1998] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (334 < i_size && h_count >= i_worm_x[2009:2004] * PIXEL_SIZE && h_count < i_worm_x[2009:2004] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2009:2004] * PIXEL_SIZE && v_count < i_worm_y[2009:2004] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (335 < i_size && h_count >= i_worm_x[2015:2010] * PIXEL_SIZE && h_count < i_worm_x[2015:2010] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2015:2010] * PIXEL_SIZE && v_count < i_worm_y[2015:2010] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (336 < i_size && h_count >= i_worm_x[2021:2016] * PIXEL_SIZE && h_count < i_worm_x[2021:2016] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2021:2016] * PIXEL_SIZE && v_count < i_worm_y[2021:2016] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (337 < i_size && h_count >= i_worm_x[2027:2022] * PIXEL_SIZE && h_count < i_worm_x[2027:2022] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2027:2022] * PIXEL_SIZE && v_count < i_worm_y[2027:2022] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (338 < i_size && h_count >= i_worm_x[2033:2028] * PIXEL_SIZE && h_count < i_worm_x[2033:2028] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2033:2028] * PIXEL_SIZE && v_count < i_worm_y[2033:2028] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (339 < i_size && h_count >= i_worm_x[2039:2034] * PIXEL_SIZE && h_count < i_worm_x[2039:2034] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2039:2034] * PIXEL_SIZE && v_count < i_worm_y[2039:2034] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (340 < i_size && h_count >= i_worm_x[2045:2040] * PIXEL_SIZE && h_count < i_worm_x[2045:2040] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2045:2040] * PIXEL_SIZE && v_count < i_worm_y[2045:2040] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (341 < i_size && h_count >= i_worm_x[2051:2046] * PIXEL_SIZE && h_count < i_worm_x[2051:2046] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2051:2046] * PIXEL_SIZE && v_count < i_worm_y[2051:2046] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (342 < i_size && h_count >= i_worm_x[2057:2052] * PIXEL_SIZE && h_count < i_worm_x[2057:2052] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2057:2052] * PIXEL_SIZE && v_count < i_worm_y[2057:2052] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (343 < i_size && h_count >= i_worm_x[2063:2058] * PIXEL_SIZE && h_count < i_worm_x[2063:2058] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2063:2058] * PIXEL_SIZE && v_count < i_worm_y[2063:2058] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (344 < i_size && h_count >= i_worm_x[2069:2064] * PIXEL_SIZE && h_count < i_worm_x[2069:2064] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2069:2064] * PIXEL_SIZE && v_count < i_worm_y[2069:2064] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (345 < i_size && h_count >= i_worm_x[2075:2070] * PIXEL_SIZE && h_count < i_worm_x[2075:2070] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2075:2070] * PIXEL_SIZE && v_count < i_worm_y[2075:2070] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (346 < i_size && h_count >= i_worm_x[2081:2076] * PIXEL_SIZE && h_count < i_worm_x[2081:2076] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2081:2076] * PIXEL_SIZE && v_count < i_worm_y[2081:2076] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (347 < i_size && h_count >= i_worm_x[2087:2082] * PIXEL_SIZE && h_count < i_worm_x[2087:2082] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2087:2082] * PIXEL_SIZE && v_count < i_worm_y[2087:2082] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (348 < i_size && h_count >= i_worm_x[2093:2088] * PIXEL_SIZE && h_count < i_worm_x[2093:2088] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2093:2088] * PIXEL_SIZE && v_count < i_worm_y[2093:2088] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (349 < i_size && h_count >= i_worm_x[2099:2094] * PIXEL_SIZE && h_count < i_worm_x[2099:2094] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2099:2094] * PIXEL_SIZE && v_count < i_worm_y[2099:2094] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (350 < i_size && h_count >= i_worm_x[2105:2100] * PIXEL_SIZE && h_count < i_worm_x[2105:2100] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2105:2100] * PIXEL_SIZE && v_count < i_worm_y[2105:2100] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (351 < i_size && h_count >= i_worm_x[2111:2106] * PIXEL_SIZE && h_count < i_worm_x[2111:2106] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2111:2106] * PIXEL_SIZE && v_count < i_worm_y[2111:2106] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (352 < i_size && h_count >= i_worm_x[2117:2112] * PIXEL_SIZE && h_count < i_worm_x[2117:2112] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2117:2112] * PIXEL_SIZE && v_count < i_worm_y[2117:2112] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (353 < i_size && h_count >= i_worm_x[2123:2118] * PIXEL_SIZE && h_count < i_worm_x[2123:2118] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2123:2118] * PIXEL_SIZE && v_count < i_worm_y[2123:2118] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (354 < i_size && h_count >= i_worm_x[2129:2124] * PIXEL_SIZE && h_count < i_worm_x[2129:2124] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2129:2124] * PIXEL_SIZE && v_count < i_worm_y[2129:2124] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (355 < i_size && h_count >= i_worm_x[2135:2130] * PIXEL_SIZE && h_count < i_worm_x[2135:2130] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2135:2130] * PIXEL_SIZE && v_count < i_worm_y[2135:2130] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (356 < i_size && h_count >= i_worm_x[2141:2136] * PIXEL_SIZE && h_count < i_worm_x[2141:2136] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2141:2136] * PIXEL_SIZE && v_count < i_worm_y[2141:2136] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (357 < i_size && h_count >= i_worm_x[2147:2142] * PIXEL_SIZE && h_count < i_worm_x[2147:2142] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2147:2142] * PIXEL_SIZE && v_count < i_worm_y[2147:2142] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (358 < i_size && h_count >= i_worm_x[2153:2148] * PIXEL_SIZE && h_count < i_worm_x[2153:2148] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2153:2148] * PIXEL_SIZE && v_count < i_worm_y[2153:2148] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (359 < i_size && h_count >= i_worm_x[2159:2154] * PIXEL_SIZE && h_count < i_worm_x[2159:2154] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2159:2154] * PIXEL_SIZE && v_count < i_worm_y[2159:2154] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (360 < i_size && h_count >= i_worm_x[2165:2160] * PIXEL_SIZE && h_count < i_worm_x[2165:2160] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2165:2160] * PIXEL_SIZE && v_count < i_worm_y[2165:2160] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (361 < i_size && h_count >= i_worm_x[2171:2166] * PIXEL_SIZE && h_count < i_worm_x[2171:2166] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2171:2166] * PIXEL_SIZE && v_count < i_worm_y[2171:2166] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (362 < i_size && h_count >= i_worm_x[2177:2172] * PIXEL_SIZE && h_count < i_worm_x[2177:2172] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2177:2172] * PIXEL_SIZE && v_count < i_worm_y[2177:2172] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (363 < i_size && h_count >= i_worm_x[2183:2178] * PIXEL_SIZE && h_count < i_worm_x[2183:2178] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2183:2178] * PIXEL_SIZE && v_count < i_worm_y[2183:2178] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (364 < i_size && h_count >= i_worm_x[2189:2184] * PIXEL_SIZE && h_count < i_worm_x[2189:2184] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2189:2184] * PIXEL_SIZE && v_count < i_worm_y[2189:2184] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (365 < i_size && h_count >= i_worm_x[2195:2190] * PIXEL_SIZE && h_count < i_worm_x[2195:2190] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2195:2190] * PIXEL_SIZE && v_count < i_worm_y[2195:2190] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (366 < i_size && h_count >= i_worm_x[2201:2196] * PIXEL_SIZE && h_count < i_worm_x[2201:2196] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2201:2196] * PIXEL_SIZE && v_count < i_worm_y[2201:2196] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (367 < i_size && h_count >= i_worm_x[2207:2202] * PIXEL_SIZE && h_count < i_worm_x[2207:2202] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2207:2202] * PIXEL_SIZE && v_count < i_worm_y[2207:2202] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (368 < i_size && h_count >= i_worm_x[2213:2208] * PIXEL_SIZE && h_count < i_worm_x[2213:2208] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2213:2208] * PIXEL_SIZE && v_count < i_worm_y[2213:2208] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (369 < i_size && h_count >= i_worm_x[2219:2214] * PIXEL_SIZE && h_count < i_worm_x[2219:2214] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2219:2214] * PIXEL_SIZE && v_count < i_worm_y[2219:2214] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (370 < i_size && h_count >= i_worm_x[2225:2220] * PIXEL_SIZE && h_count < i_worm_x[2225:2220] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2225:2220] * PIXEL_SIZE && v_count < i_worm_y[2225:2220] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (371 < i_size && h_count >= i_worm_x[2231:2226] * PIXEL_SIZE && h_count < i_worm_x[2231:2226] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2231:2226] * PIXEL_SIZE && v_count < i_worm_y[2231:2226] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (372 < i_size && h_count >= i_worm_x[2237:2232] * PIXEL_SIZE && h_count < i_worm_x[2237:2232] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2237:2232] * PIXEL_SIZE && v_count < i_worm_y[2237:2232] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (373 < i_size && h_count >= i_worm_x[2243:2238] * PIXEL_SIZE && h_count < i_worm_x[2243:2238] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2243:2238] * PIXEL_SIZE && v_count < i_worm_y[2243:2238] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (374 < i_size && h_count >= i_worm_x[2249:2244] * PIXEL_SIZE && h_count < i_worm_x[2249:2244] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2249:2244] * PIXEL_SIZE && v_count < i_worm_y[2249:2244] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (375 < i_size && h_count >= i_worm_x[2255:2250] * PIXEL_SIZE && h_count < i_worm_x[2255:2250] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2255:2250] * PIXEL_SIZE && v_count < i_worm_y[2255:2250] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (376 < i_size && h_count >= i_worm_x[2261:2256] * PIXEL_SIZE && h_count < i_worm_x[2261:2256] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2261:2256] * PIXEL_SIZE && v_count < i_worm_y[2261:2256] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (377 < i_size && h_count >= i_worm_x[2267:2262] * PIXEL_SIZE && h_count < i_worm_x[2267:2262] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2267:2262] * PIXEL_SIZE && v_count < i_worm_y[2267:2262] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (378 < i_size && h_count >= i_worm_x[2273:2268] * PIXEL_SIZE && h_count < i_worm_x[2273:2268] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2273:2268] * PIXEL_SIZE && v_count < i_worm_y[2273:2268] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (379 < i_size && h_count >= i_worm_x[2279:2274] * PIXEL_SIZE && h_count < i_worm_x[2279:2274] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2279:2274] * PIXEL_SIZE && v_count < i_worm_y[2279:2274] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (380 < i_size && h_count >= i_worm_x[2285:2280] * PIXEL_SIZE && h_count < i_worm_x[2285:2280] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2285:2280] * PIXEL_SIZE && v_count < i_worm_y[2285:2280] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (381 < i_size && h_count >= i_worm_x[2291:2286] * PIXEL_SIZE && h_count < i_worm_x[2291:2286] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2291:2286] * PIXEL_SIZE && v_count < i_worm_y[2291:2286] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (382 < i_size && h_count >= i_worm_x[2297:2292] * PIXEL_SIZE && h_count < i_worm_x[2297:2292] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2297:2292] * PIXEL_SIZE && v_count < i_worm_y[2297:2292] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (383 < i_size && h_count >= i_worm_x[2303:2298] * PIXEL_SIZE && h_count < i_worm_x[2303:2298] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2303:2298] * PIXEL_SIZE && v_count < i_worm_y[2303:2298] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (384 < i_size && h_count >= i_worm_x[2309:2304] * PIXEL_SIZE && h_count < i_worm_x[2309:2304] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2309:2304] * PIXEL_SIZE && v_count < i_worm_y[2309:2304] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (385 < i_size && h_count >= i_worm_x[2315:2310] * PIXEL_SIZE && h_count < i_worm_x[2315:2310] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2315:2310] * PIXEL_SIZE && v_count < i_worm_y[2315:2310] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (386 < i_size && h_count >= i_worm_x[2321:2316] * PIXEL_SIZE && h_count < i_worm_x[2321:2316] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2321:2316] * PIXEL_SIZE && v_count < i_worm_y[2321:2316] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (387 < i_size && h_count >= i_worm_x[2327:2322] * PIXEL_SIZE && h_count < i_worm_x[2327:2322] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2327:2322] * PIXEL_SIZE && v_count < i_worm_y[2327:2322] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (388 < i_size && h_count >= i_worm_x[2333:2328] * PIXEL_SIZE && h_count < i_worm_x[2333:2328] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2333:2328] * PIXEL_SIZE && v_count < i_worm_y[2333:2328] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (389 < i_size && h_count >= i_worm_x[2339:2334] * PIXEL_SIZE && h_count < i_worm_x[2339:2334] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2339:2334] * PIXEL_SIZE && v_count < i_worm_y[2339:2334] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (390 < i_size && h_count >= i_worm_x[2345:2340] * PIXEL_SIZE && h_count < i_worm_x[2345:2340] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2345:2340] * PIXEL_SIZE && v_count < i_worm_y[2345:2340] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (391 < i_size && h_count >= i_worm_x[2351:2346] * PIXEL_SIZE && h_count < i_worm_x[2351:2346] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2351:2346] * PIXEL_SIZE && v_count < i_worm_y[2351:2346] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (392 < i_size && h_count >= i_worm_x[2357:2352] * PIXEL_SIZE && h_count < i_worm_x[2357:2352] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2357:2352] * PIXEL_SIZE && v_count < i_worm_y[2357:2352] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (393 < i_size && h_count >= i_worm_x[2363:2358] * PIXEL_SIZE && h_count < i_worm_x[2363:2358] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2363:2358] * PIXEL_SIZE && v_count < i_worm_y[2363:2358] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (394 < i_size && h_count >= i_worm_x[2369:2364] * PIXEL_SIZE && h_count < i_worm_x[2369:2364] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2369:2364] * PIXEL_SIZE && v_count < i_worm_y[2369:2364] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (395 < i_size && h_count >= i_worm_x[2375:2370] * PIXEL_SIZE && h_count < i_worm_x[2375:2370] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2375:2370] * PIXEL_SIZE && v_count < i_worm_y[2375:2370] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (396 < i_size && h_count >= i_worm_x[2381:2376] * PIXEL_SIZE && h_count < i_worm_x[2381:2376] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2381:2376] * PIXEL_SIZE && v_count < i_worm_y[2381:2376] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (397 < i_size && h_count >= i_worm_x[2387:2382] * PIXEL_SIZE && h_count < i_worm_x[2387:2382] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2387:2382] * PIXEL_SIZE && v_count < i_worm_y[2387:2382] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (398 < i_size && h_count >= i_worm_x[2393:2388] * PIXEL_SIZE && h_count < i_worm_x[2393:2388] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2393:2388] * PIXEL_SIZE && v_count < i_worm_y[2393:2388] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (399 < i_size && h_count >= i_worm_x[2399:2394] * PIXEL_SIZE && h_count < i_worm_x[2399:2394] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2399:2394] * PIXEL_SIZE && v_count < i_worm_y[2399:2394] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (400 < i_size && h_count >= i_worm_x[2405:2400] * PIXEL_SIZE && h_count < i_worm_x[2405:2400] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2405:2400] * PIXEL_SIZE && v_count < i_worm_y[2405:2400] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (401 < i_size && h_count >= i_worm_x[2411:2406] * PIXEL_SIZE && h_count < i_worm_x[2411:2406] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2411:2406] * PIXEL_SIZE && v_count < i_worm_y[2411:2406] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (402 < i_size && h_count >= i_worm_x[2417:2412] * PIXEL_SIZE && h_count < i_worm_x[2417:2412] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2417:2412] * PIXEL_SIZE && v_count < i_worm_y[2417:2412] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (403 < i_size && h_count >= i_worm_x[2423:2418] * PIXEL_SIZE && h_count < i_worm_x[2423:2418] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2423:2418] * PIXEL_SIZE && v_count < i_worm_y[2423:2418] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (404 < i_size && h_count >= i_worm_x[2429:2424] * PIXEL_SIZE && h_count < i_worm_x[2429:2424] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2429:2424] * PIXEL_SIZE && v_count < i_worm_y[2429:2424] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (405 < i_size && h_count >= i_worm_x[2435:2430] * PIXEL_SIZE && h_count < i_worm_x[2435:2430] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2435:2430] * PIXEL_SIZE && v_count < i_worm_y[2435:2430] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (406 < i_size && h_count >= i_worm_x[2441:2436] * PIXEL_SIZE && h_count < i_worm_x[2441:2436] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2441:2436] * PIXEL_SIZE && v_count < i_worm_y[2441:2436] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (407 < i_size && h_count >= i_worm_x[2447:2442] * PIXEL_SIZE && h_count < i_worm_x[2447:2442] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2447:2442] * PIXEL_SIZE && v_count < i_worm_y[2447:2442] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (408 < i_size && h_count >= i_worm_x[2453:2448] * PIXEL_SIZE && h_count < i_worm_x[2453:2448] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2453:2448] * PIXEL_SIZE && v_count < i_worm_y[2453:2448] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (409 < i_size && h_count >= i_worm_x[2459:2454] * PIXEL_SIZE && h_count < i_worm_x[2459:2454] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2459:2454] * PIXEL_SIZE && v_count < i_worm_y[2459:2454] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (410 < i_size && h_count >= i_worm_x[2465:2460] * PIXEL_SIZE && h_count < i_worm_x[2465:2460] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2465:2460] * PIXEL_SIZE && v_count < i_worm_y[2465:2460] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (411 < i_size && h_count >= i_worm_x[2471:2466] * PIXEL_SIZE && h_count < i_worm_x[2471:2466] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2471:2466] * PIXEL_SIZE && v_count < i_worm_y[2471:2466] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (412 < i_size && h_count >= i_worm_x[2477:2472] * PIXEL_SIZE && h_count < i_worm_x[2477:2472] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2477:2472] * PIXEL_SIZE && v_count < i_worm_y[2477:2472] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (413 < i_size && h_count >= i_worm_x[2483:2478] * PIXEL_SIZE && h_count < i_worm_x[2483:2478] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2483:2478] * PIXEL_SIZE && v_count < i_worm_y[2483:2478] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (414 < i_size && h_count >= i_worm_x[2489:2484] * PIXEL_SIZE && h_count < i_worm_x[2489:2484] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2489:2484] * PIXEL_SIZE && v_count < i_worm_y[2489:2484] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (415 < i_size && h_count >= i_worm_x[2495:2490] * PIXEL_SIZE && h_count < i_worm_x[2495:2490] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2495:2490] * PIXEL_SIZE && v_count < i_worm_y[2495:2490] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (416 < i_size && h_count >= i_worm_x[2501:2496] * PIXEL_SIZE && h_count < i_worm_x[2501:2496] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2501:2496] * PIXEL_SIZE && v_count < i_worm_y[2501:2496] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (417 < i_size && h_count >= i_worm_x[2507:2502] * PIXEL_SIZE && h_count < i_worm_x[2507:2502] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2507:2502] * PIXEL_SIZE && v_count < i_worm_y[2507:2502] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (418 < i_size && h_count >= i_worm_x[2513:2508] * PIXEL_SIZE && h_count < i_worm_x[2513:2508] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2513:2508] * PIXEL_SIZE && v_count < i_worm_y[2513:2508] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (419 < i_size && h_count >= i_worm_x[2519:2514] * PIXEL_SIZE && h_count < i_worm_x[2519:2514] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2519:2514] * PIXEL_SIZE && v_count < i_worm_y[2519:2514] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (420 < i_size && h_count >= i_worm_x[2525:2520] * PIXEL_SIZE && h_count < i_worm_x[2525:2520] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2525:2520] * PIXEL_SIZE && v_count < i_worm_y[2525:2520] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (421 < i_size && h_count >= i_worm_x[2531:2526] * PIXEL_SIZE && h_count < i_worm_x[2531:2526] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2531:2526] * PIXEL_SIZE && v_count < i_worm_y[2531:2526] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (422 < i_size && h_count >= i_worm_x[2537:2532] * PIXEL_SIZE && h_count < i_worm_x[2537:2532] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2537:2532] * PIXEL_SIZE && v_count < i_worm_y[2537:2532] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (423 < i_size && h_count >= i_worm_x[2543:2538] * PIXEL_SIZE && h_count < i_worm_x[2543:2538] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2543:2538] * PIXEL_SIZE && v_count < i_worm_y[2543:2538] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (424 < i_size && h_count >= i_worm_x[2549:2544] * PIXEL_SIZE && h_count < i_worm_x[2549:2544] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2549:2544] * PIXEL_SIZE && v_count < i_worm_y[2549:2544] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (425 < i_size && h_count >= i_worm_x[2555:2550] * PIXEL_SIZE && h_count < i_worm_x[2555:2550] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2555:2550] * PIXEL_SIZE && v_count < i_worm_y[2555:2550] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (426 < i_size && h_count >= i_worm_x[2561:2556] * PIXEL_SIZE && h_count < i_worm_x[2561:2556] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2561:2556] * PIXEL_SIZE && v_count < i_worm_y[2561:2556] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (427 < i_size && h_count >= i_worm_x[2567:2562] * PIXEL_SIZE && h_count < i_worm_x[2567:2562] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2567:2562] * PIXEL_SIZE && v_count < i_worm_y[2567:2562] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (428 < i_size && h_count >= i_worm_x[2573:2568] * PIXEL_SIZE && h_count < i_worm_x[2573:2568] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2573:2568] * PIXEL_SIZE && v_count < i_worm_y[2573:2568] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (429 < i_size && h_count >= i_worm_x[2579:2574] * PIXEL_SIZE && h_count < i_worm_x[2579:2574] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2579:2574] * PIXEL_SIZE && v_count < i_worm_y[2579:2574] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (430 < i_size && h_count >= i_worm_x[2585:2580] * PIXEL_SIZE && h_count < i_worm_x[2585:2580] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2585:2580] * PIXEL_SIZE && v_count < i_worm_y[2585:2580] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (431 < i_size && h_count >= i_worm_x[2591:2586] * PIXEL_SIZE && h_count < i_worm_x[2591:2586] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2591:2586] * PIXEL_SIZE && v_count < i_worm_y[2591:2586] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (432 < i_size && h_count >= i_worm_x[2597:2592] * PIXEL_SIZE && h_count < i_worm_x[2597:2592] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2597:2592] * PIXEL_SIZE && v_count < i_worm_y[2597:2592] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (433 < i_size && h_count >= i_worm_x[2603:2598] * PIXEL_SIZE && h_count < i_worm_x[2603:2598] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2603:2598] * PIXEL_SIZE && v_count < i_worm_y[2603:2598] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (434 < i_size && h_count >= i_worm_x[2609:2604] * PIXEL_SIZE && h_count < i_worm_x[2609:2604] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2609:2604] * PIXEL_SIZE && v_count < i_worm_y[2609:2604] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (435 < i_size && h_count >= i_worm_x[2615:2610] * PIXEL_SIZE && h_count < i_worm_x[2615:2610] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2615:2610] * PIXEL_SIZE && v_count < i_worm_y[2615:2610] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (436 < i_size && h_count >= i_worm_x[2621:2616] * PIXEL_SIZE && h_count < i_worm_x[2621:2616] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2621:2616] * PIXEL_SIZE && v_count < i_worm_y[2621:2616] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (437 < i_size && h_count >= i_worm_x[2627:2622] * PIXEL_SIZE && h_count < i_worm_x[2627:2622] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2627:2622] * PIXEL_SIZE && v_count < i_worm_y[2627:2622] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (438 < i_size && h_count >= i_worm_x[2633:2628] * PIXEL_SIZE && h_count < i_worm_x[2633:2628] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2633:2628] * PIXEL_SIZE && v_count < i_worm_y[2633:2628] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (439 < i_size && h_count >= i_worm_x[2639:2634] * PIXEL_SIZE && h_count < i_worm_x[2639:2634] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2639:2634] * PIXEL_SIZE && v_count < i_worm_y[2639:2634] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (440 < i_size && h_count >= i_worm_x[2645:2640] * PIXEL_SIZE && h_count < i_worm_x[2645:2640] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2645:2640] * PIXEL_SIZE && v_count < i_worm_y[2645:2640] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (441 < i_size && h_count >= i_worm_x[2651:2646] * PIXEL_SIZE && h_count < i_worm_x[2651:2646] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2651:2646] * PIXEL_SIZE && v_count < i_worm_y[2651:2646] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (442 < i_size && h_count >= i_worm_x[2657:2652] * PIXEL_SIZE && h_count < i_worm_x[2657:2652] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2657:2652] * PIXEL_SIZE && v_count < i_worm_y[2657:2652] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (443 < i_size && h_count >= i_worm_x[2663:2658] * PIXEL_SIZE && h_count < i_worm_x[2663:2658] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2663:2658] * PIXEL_SIZE && v_count < i_worm_y[2663:2658] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (444 < i_size && h_count >= i_worm_x[2669:2664] * PIXEL_SIZE && h_count < i_worm_x[2669:2664] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2669:2664] * PIXEL_SIZE && v_count < i_worm_y[2669:2664] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (445 < i_size && h_count >= i_worm_x[2675:2670] * PIXEL_SIZE && h_count < i_worm_x[2675:2670] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2675:2670] * PIXEL_SIZE && v_count < i_worm_y[2675:2670] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (446 < i_size && h_count >= i_worm_x[2681:2676] * PIXEL_SIZE && h_count < i_worm_x[2681:2676] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2681:2676] * PIXEL_SIZE && v_count < i_worm_y[2681:2676] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (447 < i_size && h_count >= i_worm_x[2687:2682] * PIXEL_SIZE && h_count < i_worm_x[2687:2682] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2687:2682] * PIXEL_SIZE && v_count < i_worm_y[2687:2682] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (448 < i_size && h_count >= i_worm_x[2693:2688] * PIXEL_SIZE && h_count < i_worm_x[2693:2688] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2693:2688] * PIXEL_SIZE && v_count < i_worm_y[2693:2688] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (449 < i_size && h_count >= i_worm_x[2699:2694] * PIXEL_SIZE && h_count < i_worm_x[2699:2694] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2699:2694] * PIXEL_SIZE && v_count < i_worm_y[2699:2694] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (450 < i_size && h_count >= i_worm_x[2705:2700] * PIXEL_SIZE && h_count < i_worm_x[2705:2700] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2705:2700] * PIXEL_SIZE && v_count < i_worm_y[2705:2700] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (451 < i_size && h_count >= i_worm_x[2711:2706] * PIXEL_SIZE && h_count < i_worm_x[2711:2706] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2711:2706] * PIXEL_SIZE && v_count < i_worm_y[2711:2706] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (452 < i_size && h_count >= i_worm_x[2717:2712] * PIXEL_SIZE && h_count < i_worm_x[2717:2712] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2717:2712] * PIXEL_SIZE && v_count < i_worm_y[2717:2712] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (453 < i_size && h_count >= i_worm_x[2723:2718] * PIXEL_SIZE && h_count < i_worm_x[2723:2718] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2723:2718] * PIXEL_SIZE && v_count < i_worm_y[2723:2718] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (454 < i_size && h_count >= i_worm_x[2729:2724] * PIXEL_SIZE && h_count < i_worm_x[2729:2724] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2729:2724] * PIXEL_SIZE && v_count < i_worm_y[2729:2724] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (455 < i_size && h_count >= i_worm_x[2735:2730] * PIXEL_SIZE && h_count < i_worm_x[2735:2730] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2735:2730] * PIXEL_SIZE && v_count < i_worm_y[2735:2730] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (456 < i_size && h_count >= i_worm_x[2741:2736] * PIXEL_SIZE && h_count < i_worm_x[2741:2736] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2741:2736] * PIXEL_SIZE && v_count < i_worm_y[2741:2736] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (457 < i_size && h_count >= i_worm_x[2747:2742] * PIXEL_SIZE && h_count < i_worm_x[2747:2742] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2747:2742] * PIXEL_SIZE && v_count < i_worm_y[2747:2742] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (458 < i_size && h_count >= i_worm_x[2753:2748] * PIXEL_SIZE && h_count < i_worm_x[2753:2748] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2753:2748] * PIXEL_SIZE && v_count < i_worm_y[2753:2748] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (459 < i_size && h_count >= i_worm_x[2759:2754] * PIXEL_SIZE && h_count < i_worm_x[2759:2754] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2759:2754] * PIXEL_SIZE && v_count < i_worm_y[2759:2754] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (460 < i_size && h_count >= i_worm_x[2765:2760] * PIXEL_SIZE && h_count < i_worm_x[2765:2760] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2765:2760] * PIXEL_SIZE && v_count < i_worm_y[2765:2760] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (461 < i_size && h_count >= i_worm_x[2771:2766] * PIXEL_SIZE && h_count < i_worm_x[2771:2766] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2771:2766] * PIXEL_SIZE && v_count < i_worm_y[2771:2766] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (462 < i_size && h_count >= i_worm_x[2777:2772] * PIXEL_SIZE && h_count < i_worm_x[2777:2772] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2777:2772] * PIXEL_SIZE && v_count < i_worm_y[2777:2772] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (463 < i_size && h_count >= i_worm_x[2783:2778] * PIXEL_SIZE && h_count < i_worm_x[2783:2778] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2783:2778] * PIXEL_SIZE && v_count < i_worm_y[2783:2778] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (464 < i_size && h_count >= i_worm_x[2789:2784] * PIXEL_SIZE && h_count < i_worm_x[2789:2784] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2789:2784] * PIXEL_SIZE && v_count < i_worm_y[2789:2784] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (465 < i_size && h_count >= i_worm_x[2795:2790] * PIXEL_SIZE && h_count < i_worm_x[2795:2790] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2795:2790] * PIXEL_SIZE && v_count < i_worm_y[2795:2790] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (466 < i_size && h_count >= i_worm_x[2801:2796] * PIXEL_SIZE && h_count < i_worm_x[2801:2796] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2801:2796] * PIXEL_SIZE && v_count < i_worm_y[2801:2796] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (467 < i_size && h_count >= i_worm_x[2807:2802] * PIXEL_SIZE && h_count < i_worm_x[2807:2802] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2807:2802] * PIXEL_SIZE && v_count < i_worm_y[2807:2802] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (468 < i_size && h_count >= i_worm_x[2813:2808] * PIXEL_SIZE && h_count < i_worm_x[2813:2808] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2813:2808] * PIXEL_SIZE && v_count < i_worm_y[2813:2808] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (469 < i_size && h_count >= i_worm_x[2819:2814] * PIXEL_SIZE && h_count < i_worm_x[2819:2814] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2819:2814] * PIXEL_SIZE && v_count < i_worm_y[2819:2814] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (470 < i_size && h_count >= i_worm_x[2825:2820] * PIXEL_SIZE && h_count < i_worm_x[2825:2820] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2825:2820] * PIXEL_SIZE && v_count < i_worm_y[2825:2820] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (471 < i_size && h_count >= i_worm_x[2831:2826] * PIXEL_SIZE && h_count < i_worm_x[2831:2826] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2831:2826] * PIXEL_SIZE && v_count < i_worm_y[2831:2826] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (472 < i_size && h_count >= i_worm_x[2837:2832] * PIXEL_SIZE && h_count < i_worm_x[2837:2832] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2837:2832] * PIXEL_SIZE && v_count < i_worm_y[2837:2832] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (473 < i_size && h_count >= i_worm_x[2843:2838] * PIXEL_SIZE && h_count < i_worm_x[2843:2838] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2843:2838] * PIXEL_SIZE && v_count < i_worm_y[2843:2838] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (474 < i_size && h_count >= i_worm_x[2849:2844] * PIXEL_SIZE && h_count < i_worm_x[2849:2844] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2849:2844] * PIXEL_SIZE && v_count < i_worm_y[2849:2844] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (475 < i_size && h_count >= i_worm_x[2855:2850] * PIXEL_SIZE && h_count < i_worm_x[2855:2850] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2855:2850] * PIXEL_SIZE && v_count < i_worm_y[2855:2850] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (476 < i_size && h_count >= i_worm_x[2861:2856] * PIXEL_SIZE && h_count < i_worm_x[2861:2856] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2861:2856] * PIXEL_SIZE && v_count < i_worm_y[2861:2856] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (477 < i_size && h_count >= i_worm_x[2867:2862] * PIXEL_SIZE && h_count < i_worm_x[2867:2862] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2867:2862] * PIXEL_SIZE && v_count < i_worm_y[2867:2862] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (478 < i_size && h_count >= i_worm_x[2873:2868] * PIXEL_SIZE && h_count < i_worm_x[2873:2868] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2873:2868] * PIXEL_SIZE && v_count < i_worm_y[2873:2868] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (479 < i_size && h_count >= i_worm_x[2879:2874] * PIXEL_SIZE && h_count < i_worm_x[2879:2874] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2879:2874] * PIXEL_SIZE && v_count < i_worm_y[2879:2874] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (480 < i_size && h_count >= i_worm_x[2885:2880] * PIXEL_SIZE && h_count < i_worm_x[2885:2880] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2885:2880] * PIXEL_SIZE && v_count < i_worm_y[2885:2880] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (481 < i_size && h_count >= i_worm_x[2891:2886] * PIXEL_SIZE && h_count < i_worm_x[2891:2886] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2891:2886] * PIXEL_SIZE && v_count < i_worm_y[2891:2886] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (482 < i_size && h_count >= i_worm_x[2897:2892] * PIXEL_SIZE && h_count < i_worm_x[2897:2892] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2897:2892] * PIXEL_SIZE && v_count < i_worm_y[2897:2892] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (483 < i_size && h_count >= i_worm_x[2903:2898] * PIXEL_SIZE && h_count < i_worm_x[2903:2898] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2903:2898] * PIXEL_SIZE && v_count < i_worm_y[2903:2898] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (484 < i_size && h_count >= i_worm_x[2909:2904] * PIXEL_SIZE && h_count < i_worm_x[2909:2904] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2909:2904] * PIXEL_SIZE && v_count < i_worm_y[2909:2904] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (485 < i_size && h_count >= i_worm_x[2915:2910] * PIXEL_SIZE && h_count < i_worm_x[2915:2910] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2915:2910] * PIXEL_SIZE && v_count < i_worm_y[2915:2910] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (486 < i_size && h_count >= i_worm_x[2921:2916] * PIXEL_SIZE && h_count < i_worm_x[2921:2916] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2921:2916] * PIXEL_SIZE && v_count < i_worm_y[2921:2916] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (487 < i_size && h_count >= i_worm_x[2927:2922] * PIXEL_SIZE && h_count < i_worm_x[2927:2922] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2927:2922] * PIXEL_SIZE && v_count < i_worm_y[2927:2922] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (488 < i_size && h_count >= i_worm_x[2933:2928] * PIXEL_SIZE && h_count < i_worm_x[2933:2928] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2933:2928] * PIXEL_SIZE && v_count < i_worm_y[2933:2928] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (489 < i_size && h_count >= i_worm_x[2939:2934] * PIXEL_SIZE && h_count < i_worm_x[2939:2934] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2939:2934] * PIXEL_SIZE && v_count < i_worm_y[2939:2934] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (490 < i_size && h_count >= i_worm_x[2945:2940] * PIXEL_SIZE && h_count < i_worm_x[2945:2940] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2945:2940] * PIXEL_SIZE && v_count < i_worm_y[2945:2940] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (491 < i_size && h_count >= i_worm_x[2951:2946] * PIXEL_SIZE && h_count < i_worm_x[2951:2946] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2951:2946] * PIXEL_SIZE && v_count < i_worm_y[2951:2946] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (492 < i_size && h_count >= i_worm_x[2957:2952] * PIXEL_SIZE && h_count < i_worm_x[2957:2952] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2957:2952] * PIXEL_SIZE && v_count < i_worm_y[2957:2952] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (493 < i_size && h_count >= i_worm_x[2963:2958] * PIXEL_SIZE && h_count < i_worm_x[2963:2958] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2963:2958] * PIXEL_SIZE && v_count < i_worm_y[2963:2958] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (494 < i_size && h_count >= i_worm_x[2969:2964] * PIXEL_SIZE && h_count < i_worm_x[2969:2964] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2969:2964] * PIXEL_SIZE && v_count < i_worm_y[2969:2964] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (495 < i_size && h_count >= i_worm_x[2975:2970] * PIXEL_SIZE && h_count < i_worm_x[2975:2970] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2975:2970] * PIXEL_SIZE && v_count < i_worm_y[2975:2970] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (496 < i_size && h_count >= i_worm_x[2981:2976] * PIXEL_SIZE && h_count < i_worm_x[2981:2976] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2981:2976] * PIXEL_SIZE && v_count < i_worm_y[2981:2976] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (497 < i_size && h_count >= i_worm_x[2987:2982] * PIXEL_SIZE && h_count < i_worm_x[2987:2982] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2987:2982] * PIXEL_SIZE && v_count < i_worm_y[2987:2982] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (498 < i_size && h_count >= i_worm_x[2993:2988] * PIXEL_SIZE && h_count < i_worm_x[2993:2988] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2993:2988] * PIXEL_SIZE && v_count < i_worm_y[2993:2988] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (499 < i_size && h_count >= i_worm_x[2999:2994] * PIXEL_SIZE && h_count < i_worm_x[2999:2994] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[2999:2994] * PIXEL_SIZE && v_count < i_worm_y[2999:2994] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (500 < i_size && h_count >= i_worm_x[3005:3000] * PIXEL_SIZE && h_count < i_worm_x[3005:3000] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3005:3000] * PIXEL_SIZE && v_count < i_worm_y[3005:3000] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (501 < i_size && h_count >= i_worm_x[3011:3006] * PIXEL_SIZE && h_count < i_worm_x[3011:3006] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3011:3006] * PIXEL_SIZE && v_count < i_worm_y[3011:3006] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (502 < i_size && h_count >= i_worm_x[3017:3012] * PIXEL_SIZE && h_count < i_worm_x[3017:3012] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3017:3012] * PIXEL_SIZE && v_count < i_worm_y[3017:3012] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (503 < i_size && h_count >= i_worm_x[3023:3018] * PIXEL_SIZE && h_count < i_worm_x[3023:3018] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3023:3018] * PIXEL_SIZE && v_count < i_worm_y[3023:3018] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (504 < i_size && h_count >= i_worm_x[3029:3024] * PIXEL_SIZE && h_count < i_worm_x[3029:3024] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3029:3024] * PIXEL_SIZE && v_count < i_worm_y[3029:3024] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (505 < i_size && h_count >= i_worm_x[3035:3030] * PIXEL_SIZE && h_count < i_worm_x[3035:3030] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3035:3030] * PIXEL_SIZE && v_count < i_worm_y[3035:3030] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (506 < i_size && h_count >= i_worm_x[3041:3036] * PIXEL_SIZE && h_count < i_worm_x[3041:3036] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3041:3036] * PIXEL_SIZE && v_count < i_worm_y[3041:3036] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (507 < i_size && h_count >= i_worm_x[3047:3042] * PIXEL_SIZE && h_count < i_worm_x[3047:3042] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3047:3042] * PIXEL_SIZE && v_count < i_worm_y[3047:3042] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (508 < i_size && h_count >= i_worm_x[3053:3048] * PIXEL_SIZE && h_count < i_worm_x[3053:3048] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3053:3048] * PIXEL_SIZE && v_count < i_worm_y[3053:3048] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (509 < i_size && h_count >= i_worm_x[3059:3054] * PIXEL_SIZE && h_count < i_worm_x[3059:3054] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3059:3054] * PIXEL_SIZE && v_count < i_worm_y[3059:3054] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (510 < i_size && h_count >= i_worm_x[3065:3060] * PIXEL_SIZE && h_count < i_worm_x[3065:3060] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3065:3060] * PIXEL_SIZE && v_count < i_worm_y[3065:3060] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (511 < i_size && h_count >= i_worm_x[3071:3066] * PIXEL_SIZE && h_count < i_worm_x[3071:3066] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3071:3066] * PIXEL_SIZE && v_count < i_worm_y[3071:3066] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (512 < i_size && h_count >= i_worm_x[3077:3072] * PIXEL_SIZE && h_count < i_worm_x[3077:3072] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3077:3072] * PIXEL_SIZE && v_count < i_worm_y[3077:3072] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (513 < i_size && h_count >= i_worm_x[3083:3078] * PIXEL_SIZE && h_count < i_worm_x[3083:3078] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3083:3078] * PIXEL_SIZE && v_count < i_worm_y[3083:3078] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (514 < i_size && h_count >= i_worm_x[3089:3084] * PIXEL_SIZE && h_count < i_worm_x[3089:3084] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3089:3084] * PIXEL_SIZE && v_count < i_worm_y[3089:3084] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (515 < i_size && h_count >= i_worm_x[3095:3090] * PIXEL_SIZE && h_count < i_worm_x[3095:3090] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3095:3090] * PIXEL_SIZE && v_count < i_worm_y[3095:3090] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (516 < i_size && h_count >= i_worm_x[3101:3096] * PIXEL_SIZE && h_count < i_worm_x[3101:3096] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3101:3096] * PIXEL_SIZE && v_count < i_worm_y[3101:3096] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (517 < i_size && h_count >= i_worm_x[3107:3102] * PIXEL_SIZE && h_count < i_worm_x[3107:3102] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3107:3102] * PIXEL_SIZE && v_count < i_worm_y[3107:3102] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (518 < i_size && h_count >= i_worm_x[3113:3108] * PIXEL_SIZE && h_count < i_worm_x[3113:3108] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3113:3108] * PIXEL_SIZE && v_count < i_worm_y[3113:3108] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (519 < i_size && h_count >= i_worm_x[3119:3114] * PIXEL_SIZE && h_count < i_worm_x[3119:3114] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3119:3114] * PIXEL_SIZE && v_count < i_worm_y[3119:3114] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (520 < i_size && h_count >= i_worm_x[3125:3120] * PIXEL_SIZE && h_count < i_worm_x[3125:3120] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3125:3120] * PIXEL_SIZE && v_count < i_worm_y[3125:3120] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (521 < i_size && h_count >= i_worm_x[3131:3126] * PIXEL_SIZE && h_count < i_worm_x[3131:3126] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3131:3126] * PIXEL_SIZE && v_count < i_worm_y[3131:3126] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (522 < i_size && h_count >= i_worm_x[3137:3132] * PIXEL_SIZE && h_count < i_worm_x[3137:3132] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3137:3132] * PIXEL_SIZE && v_count < i_worm_y[3137:3132] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (523 < i_size && h_count >= i_worm_x[3143:3138] * PIXEL_SIZE && h_count < i_worm_x[3143:3138] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3143:3138] * PIXEL_SIZE && v_count < i_worm_y[3143:3138] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (524 < i_size && h_count >= i_worm_x[3149:3144] * PIXEL_SIZE && h_count < i_worm_x[3149:3144] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3149:3144] * PIXEL_SIZE && v_count < i_worm_y[3149:3144] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (525 < i_size && h_count >= i_worm_x[3155:3150] * PIXEL_SIZE && h_count < i_worm_x[3155:3150] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3155:3150] * PIXEL_SIZE && v_count < i_worm_y[3155:3150] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (526 < i_size && h_count >= i_worm_x[3161:3156] * PIXEL_SIZE && h_count < i_worm_x[3161:3156] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3161:3156] * PIXEL_SIZE && v_count < i_worm_y[3161:3156] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (527 < i_size && h_count >= i_worm_x[3167:3162] * PIXEL_SIZE && h_count < i_worm_x[3167:3162] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3167:3162] * PIXEL_SIZE && v_count < i_worm_y[3167:3162] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (528 < i_size && h_count >= i_worm_x[3173:3168] * PIXEL_SIZE && h_count < i_worm_x[3173:3168] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3173:3168] * PIXEL_SIZE && v_count < i_worm_y[3173:3168] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (529 < i_size && h_count >= i_worm_x[3179:3174] * PIXEL_SIZE && h_count < i_worm_x[3179:3174] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3179:3174] * PIXEL_SIZE && v_count < i_worm_y[3179:3174] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (530 < i_size && h_count >= i_worm_x[3185:3180] * PIXEL_SIZE && h_count < i_worm_x[3185:3180] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3185:3180] * PIXEL_SIZE && v_count < i_worm_y[3185:3180] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (531 < i_size && h_count >= i_worm_x[3191:3186] * PIXEL_SIZE && h_count < i_worm_x[3191:3186] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3191:3186] * PIXEL_SIZE && v_count < i_worm_y[3191:3186] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (532 < i_size && h_count >= i_worm_x[3197:3192] * PIXEL_SIZE && h_count < i_worm_x[3197:3192] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3197:3192] * PIXEL_SIZE && v_count < i_worm_y[3197:3192] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (533 < i_size && h_count >= i_worm_x[3203:3198] * PIXEL_SIZE && h_count < i_worm_x[3203:3198] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3203:3198] * PIXEL_SIZE && v_count < i_worm_y[3203:3198] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (534 < i_size && h_count >= i_worm_x[3209:3204] * PIXEL_SIZE && h_count < i_worm_x[3209:3204] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3209:3204] * PIXEL_SIZE && v_count < i_worm_y[3209:3204] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (535 < i_size && h_count >= i_worm_x[3215:3210] * PIXEL_SIZE && h_count < i_worm_x[3215:3210] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3215:3210] * PIXEL_SIZE && v_count < i_worm_y[3215:3210] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (536 < i_size && h_count >= i_worm_x[3221:3216] * PIXEL_SIZE && h_count < i_worm_x[3221:3216] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3221:3216] * PIXEL_SIZE && v_count < i_worm_y[3221:3216] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (537 < i_size && h_count >= i_worm_x[3227:3222] * PIXEL_SIZE && h_count < i_worm_x[3227:3222] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3227:3222] * PIXEL_SIZE && v_count < i_worm_y[3227:3222] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (538 < i_size && h_count >= i_worm_x[3233:3228] * PIXEL_SIZE && h_count < i_worm_x[3233:3228] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3233:3228] * PIXEL_SIZE && v_count < i_worm_y[3233:3228] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (539 < i_size && h_count >= i_worm_x[3239:3234] * PIXEL_SIZE && h_count < i_worm_x[3239:3234] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3239:3234] * PIXEL_SIZE && v_count < i_worm_y[3239:3234] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (540 < i_size && h_count >= i_worm_x[3245:3240] * PIXEL_SIZE && h_count < i_worm_x[3245:3240] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3245:3240] * PIXEL_SIZE && v_count < i_worm_y[3245:3240] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (541 < i_size && h_count >= i_worm_x[3251:3246] * PIXEL_SIZE && h_count < i_worm_x[3251:3246] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3251:3246] * PIXEL_SIZE && v_count < i_worm_y[3251:3246] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (542 < i_size && h_count >= i_worm_x[3257:3252] * PIXEL_SIZE && h_count < i_worm_x[3257:3252] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3257:3252] * PIXEL_SIZE && v_count < i_worm_y[3257:3252] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (543 < i_size && h_count >= i_worm_x[3263:3258] * PIXEL_SIZE && h_count < i_worm_x[3263:3258] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3263:3258] * PIXEL_SIZE && v_count < i_worm_y[3263:3258] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (544 < i_size && h_count >= i_worm_x[3269:3264] * PIXEL_SIZE && h_count < i_worm_x[3269:3264] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3269:3264] * PIXEL_SIZE && v_count < i_worm_y[3269:3264] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (545 < i_size && h_count >= i_worm_x[3275:3270] * PIXEL_SIZE && h_count < i_worm_x[3275:3270] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3275:3270] * PIXEL_SIZE && v_count < i_worm_y[3275:3270] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (546 < i_size && h_count >= i_worm_x[3281:3276] * PIXEL_SIZE && h_count < i_worm_x[3281:3276] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3281:3276] * PIXEL_SIZE && v_count < i_worm_y[3281:3276] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (547 < i_size && h_count >= i_worm_x[3287:3282] * PIXEL_SIZE && h_count < i_worm_x[3287:3282] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3287:3282] * PIXEL_SIZE && v_count < i_worm_y[3287:3282] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (548 < i_size && h_count >= i_worm_x[3293:3288] * PIXEL_SIZE && h_count < i_worm_x[3293:3288] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3293:3288] * PIXEL_SIZE && v_count < i_worm_y[3293:3288] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (549 < i_size && h_count >= i_worm_x[3299:3294] * PIXEL_SIZE && h_count < i_worm_x[3299:3294] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3299:3294] * PIXEL_SIZE && v_count < i_worm_y[3299:3294] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (550 < i_size && h_count >= i_worm_x[3305:3300] * PIXEL_SIZE && h_count < i_worm_x[3305:3300] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3305:3300] * PIXEL_SIZE && v_count < i_worm_y[3305:3300] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (551 < i_size && h_count >= i_worm_x[3311:3306] * PIXEL_SIZE && h_count < i_worm_x[3311:3306] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3311:3306] * PIXEL_SIZE && v_count < i_worm_y[3311:3306] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (552 < i_size && h_count >= i_worm_x[3317:3312] * PIXEL_SIZE && h_count < i_worm_x[3317:3312] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3317:3312] * PIXEL_SIZE && v_count < i_worm_y[3317:3312] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (553 < i_size && h_count >= i_worm_x[3323:3318] * PIXEL_SIZE && h_count < i_worm_x[3323:3318] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3323:3318] * PIXEL_SIZE && v_count < i_worm_y[3323:3318] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (554 < i_size && h_count >= i_worm_x[3329:3324] * PIXEL_SIZE && h_count < i_worm_x[3329:3324] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3329:3324] * PIXEL_SIZE && v_count < i_worm_y[3329:3324] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (555 < i_size && h_count >= i_worm_x[3335:3330] * PIXEL_SIZE && h_count < i_worm_x[3335:3330] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3335:3330] * PIXEL_SIZE && v_count < i_worm_y[3335:3330] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (556 < i_size && h_count >= i_worm_x[3341:3336] * PIXEL_SIZE && h_count < i_worm_x[3341:3336] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3341:3336] * PIXEL_SIZE && v_count < i_worm_y[3341:3336] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (557 < i_size && h_count >= i_worm_x[3347:3342] * PIXEL_SIZE && h_count < i_worm_x[3347:3342] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3347:3342] * PIXEL_SIZE && v_count < i_worm_y[3347:3342] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (558 < i_size && h_count >= i_worm_x[3353:3348] * PIXEL_SIZE && h_count < i_worm_x[3353:3348] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3353:3348] * PIXEL_SIZE && v_count < i_worm_y[3353:3348] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (559 < i_size && h_count >= i_worm_x[3359:3354] * PIXEL_SIZE && h_count < i_worm_x[3359:3354] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3359:3354] * PIXEL_SIZE && v_count < i_worm_y[3359:3354] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (560 < i_size && h_count >= i_worm_x[3365:3360] * PIXEL_SIZE && h_count < i_worm_x[3365:3360] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3365:3360] * PIXEL_SIZE && v_count < i_worm_y[3365:3360] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (561 < i_size && h_count >= i_worm_x[3371:3366] * PIXEL_SIZE && h_count < i_worm_x[3371:3366] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3371:3366] * PIXEL_SIZE && v_count < i_worm_y[3371:3366] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (562 < i_size && h_count >= i_worm_x[3377:3372] * PIXEL_SIZE && h_count < i_worm_x[3377:3372] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3377:3372] * PIXEL_SIZE && v_count < i_worm_y[3377:3372] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (563 < i_size && h_count >= i_worm_x[3383:3378] * PIXEL_SIZE && h_count < i_worm_x[3383:3378] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3383:3378] * PIXEL_SIZE && v_count < i_worm_y[3383:3378] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (564 < i_size && h_count >= i_worm_x[3389:3384] * PIXEL_SIZE && h_count < i_worm_x[3389:3384] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3389:3384] * PIXEL_SIZE && v_count < i_worm_y[3389:3384] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (565 < i_size && h_count >= i_worm_x[3395:3390] * PIXEL_SIZE && h_count < i_worm_x[3395:3390] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3395:3390] * PIXEL_SIZE && v_count < i_worm_y[3395:3390] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (566 < i_size && h_count >= i_worm_x[3401:3396] * PIXEL_SIZE && h_count < i_worm_x[3401:3396] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3401:3396] * PIXEL_SIZE && v_count < i_worm_y[3401:3396] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (567 < i_size && h_count >= i_worm_x[3407:3402] * PIXEL_SIZE && h_count < i_worm_x[3407:3402] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3407:3402] * PIXEL_SIZE && v_count < i_worm_y[3407:3402] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (568 < i_size && h_count >= i_worm_x[3413:3408] * PIXEL_SIZE && h_count < i_worm_x[3413:3408] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3413:3408] * PIXEL_SIZE && v_count < i_worm_y[3413:3408] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (569 < i_size && h_count >= i_worm_x[3419:3414] * PIXEL_SIZE && h_count < i_worm_x[3419:3414] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3419:3414] * PIXEL_SIZE && v_count < i_worm_y[3419:3414] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (570 < i_size && h_count >= i_worm_x[3425:3420] * PIXEL_SIZE && h_count < i_worm_x[3425:3420] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3425:3420] * PIXEL_SIZE && v_count < i_worm_y[3425:3420] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (571 < i_size && h_count >= i_worm_x[3431:3426] * PIXEL_SIZE && h_count < i_worm_x[3431:3426] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3431:3426] * PIXEL_SIZE && v_count < i_worm_y[3431:3426] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (572 < i_size && h_count >= i_worm_x[3437:3432] * PIXEL_SIZE && h_count < i_worm_x[3437:3432] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3437:3432] * PIXEL_SIZE && v_count < i_worm_y[3437:3432] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (573 < i_size && h_count >= i_worm_x[3443:3438] * PIXEL_SIZE && h_count < i_worm_x[3443:3438] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3443:3438] * PIXEL_SIZE && v_count < i_worm_y[3443:3438] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (574 < i_size && h_count >= i_worm_x[3449:3444] * PIXEL_SIZE && h_count < i_worm_x[3449:3444] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3449:3444] * PIXEL_SIZE && v_count < i_worm_y[3449:3444] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (575 < i_size && h_count >= i_worm_x[3455:3450] * PIXEL_SIZE && h_count < i_worm_x[3455:3450] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3455:3450] * PIXEL_SIZE && v_count < i_worm_y[3455:3450] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (576 < i_size && h_count >= i_worm_x[3461:3456] * PIXEL_SIZE && h_count < i_worm_x[3461:3456] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3461:3456] * PIXEL_SIZE && v_count < i_worm_y[3461:3456] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (577 < i_size && h_count >= i_worm_x[3467:3462] * PIXEL_SIZE && h_count < i_worm_x[3467:3462] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3467:3462] * PIXEL_SIZE && v_count < i_worm_y[3467:3462] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (578 < i_size && h_count >= i_worm_x[3473:3468] * PIXEL_SIZE && h_count < i_worm_x[3473:3468] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3473:3468] * PIXEL_SIZE && v_count < i_worm_y[3473:3468] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (579 < i_size && h_count >= i_worm_x[3479:3474] * PIXEL_SIZE && h_count < i_worm_x[3479:3474] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3479:3474] * PIXEL_SIZE && v_count < i_worm_y[3479:3474] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (580 < i_size && h_count >= i_worm_x[3485:3480] * PIXEL_SIZE && h_count < i_worm_x[3485:3480] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3485:3480] * PIXEL_SIZE && v_count < i_worm_y[3485:3480] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (581 < i_size && h_count >= i_worm_x[3491:3486] * PIXEL_SIZE && h_count < i_worm_x[3491:3486] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3491:3486] * PIXEL_SIZE && v_count < i_worm_y[3491:3486] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (582 < i_size && h_count >= i_worm_x[3497:3492] * PIXEL_SIZE && h_count < i_worm_x[3497:3492] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3497:3492] * PIXEL_SIZE && v_count < i_worm_y[3497:3492] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (583 < i_size && h_count >= i_worm_x[3503:3498] * PIXEL_SIZE && h_count < i_worm_x[3503:3498] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3503:3498] * PIXEL_SIZE && v_count < i_worm_y[3503:3498] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (584 < i_size && h_count >= i_worm_x[3509:3504] * PIXEL_SIZE && h_count < i_worm_x[3509:3504] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3509:3504] * PIXEL_SIZE && v_count < i_worm_y[3509:3504] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (585 < i_size && h_count >= i_worm_x[3515:3510] * PIXEL_SIZE && h_count < i_worm_x[3515:3510] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3515:3510] * PIXEL_SIZE && v_count < i_worm_y[3515:3510] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (586 < i_size && h_count >= i_worm_x[3521:3516] * PIXEL_SIZE && h_count < i_worm_x[3521:3516] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3521:3516] * PIXEL_SIZE && v_count < i_worm_y[3521:3516] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (587 < i_size && h_count >= i_worm_x[3527:3522] * PIXEL_SIZE && h_count < i_worm_x[3527:3522] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3527:3522] * PIXEL_SIZE && v_count < i_worm_y[3527:3522] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (588 < i_size && h_count >= i_worm_x[3533:3528] * PIXEL_SIZE && h_count < i_worm_x[3533:3528] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3533:3528] * PIXEL_SIZE && v_count < i_worm_y[3533:3528] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (589 < i_size && h_count >= i_worm_x[3539:3534] * PIXEL_SIZE && h_count < i_worm_x[3539:3534] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3539:3534] * PIXEL_SIZE && v_count < i_worm_y[3539:3534] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (590 < i_size && h_count >= i_worm_x[3545:3540] * PIXEL_SIZE && h_count < i_worm_x[3545:3540] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3545:3540] * PIXEL_SIZE && v_count < i_worm_y[3545:3540] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (591 < i_size && h_count >= i_worm_x[3551:3546] * PIXEL_SIZE && h_count < i_worm_x[3551:3546] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3551:3546] * PIXEL_SIZE && v_count < i_worm_y[3551:3546] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (592 < i_size && h_count >= i_worm_x[3557:3552] * PIXEL_SIZE && h_count < i_worm_x[3557:3552] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3557:3552] * PIXEL_SIZE && v_count < i_worm_y[3557:3552] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (593 < i_size && h_count >= i_worm_x[3563:3558] * PIXEL_SIZE && h_count < i_worm_x[3563:3558] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3563:3558] * PIXEL_SIZE && v_count < i_worm_y[3563:3558] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (594 < i_size && h_count >= i_worm_x[3569:3564] * PIXEL_SIZE && h_count < i_worm_x[3569:3564] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3569:3564] * PIXEL_SIZE && v_count < i_worm_y[3569:3564] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (595 < i_size && h_count >= i_worm_x[3575:3570] * PIXEL_SIZE && h_count < i_worm_x[3575:3570] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3575:3570] * PIXEL_SIZE && v_count < i_worm_y[3575:3570] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (596 < i_size && h_count >= i_worm_x[3581:3576] * PIXEL_SIZE && h_count < i_worm_x[3581:3576] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3581:3576] * PIXEL_SIZE && v_count < i_worm_y[3581:3576] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (597 < i_size && h_count >= i_worm_x[3587:3582] * PIXEL_SIZE && h_count < i_worm_x[3587:3582] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3587:3582] * PIXEL_SIZE && v_count < i_worm_y[3587:3582] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (598 < i_size && h_count >= i_worm_x[3593:3588] * PIXEL_SIZE && h_count < i_worm_x[3593:3588] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3593:3588] * PIXEL_SIZE && v_count < i_worm_y[3593:3588] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (599 < i_size && h_count >= i_worm_x[3599:3594] * PIXEL_SIZE && h_count < i_worm_x[3599:3594] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3599:3594] * PIXEL_SIZE && v_count < i_worm_y[3599:3594] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (600 < i_size && h_count >= i_worm_x[3605:3600] * PIXEL_SIZE && h_count < i_worm_x[3605:3600] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3605:3600] * PIXEL_SIZE && v_count < i_worm_y[3605:3600] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (601 < i_size && h_count >= i_worm_x[3611:3606] * PIXEL_SIZE && h_count < i_worm_x[3611:3606] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3611:3606] * PIXEL_SIZE && v_count < i_worm_y[3611:3606] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (602 < i_size && h_count >= i_worm_x[3617:3612] * PIXEL_SIZE && h_count < i_worm_x[3617:3612] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3617:3612] * PIXEL_SIZE && v_count < i_worm_y[3617:3612] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (603 < i_size && h_count >= i_worm_x[3623:3618] * PIXEL_SIZE && h_count < i_worm_x[3623:3618] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3623:3618] * PIXEL_SIZE && v_count < i_worm_y[3623:3618] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (604 < i_size && h_count >= i_worm_x[3629:3624] * PIXEL_SIZE && h_count < i_worm_x[3629:3624] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3629:3624] * PIXEL_SIZE && v_count < i_worm_y[3629:3624] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (605 < i_size && h_count >= i_worm_x[3635:3630] * PIXEL_SIZE && h_count < i_worm_x[3635:3630] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3635:3630] * PIXEL_SIZE && v_count < i_worm_y[3635:3630] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (606 < i_size && h_count >= i_worm_x[3641:3636] * PIXEL_SIZE && h_count < i_worm_x[3641:3636] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3641:3636] * PIXEL_SIZE && v_count < i_worm_y[3641:3636] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (607 < i_size && h_count >= i_worm_x[3647:3642] * PIXEL_SIZE && h_count < i_worm_x[3647:3642] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3647:3642] * PIXEL_SIZE && v_count < i_worm_y[3647:3642] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (608 < i_size && h_count >= i_worm_x[3653:3648] * PIXEL_SIZE && h_count < i_worm_x[3653:3648] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3653:3648] * PIXEL_SIZE && v_count < i_worm_y[3653:3648] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (609 < i_size && h_count >= i_worm_x[3659:3654] * PIXEL_SIZE && h_count < i_worm_x[3659:3654] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3659:3654] * PIXEL_SIZE && v_count < i_worm_y[3659:3654] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (610 < i_size && h_count >= i_worm_x[3665:3660] * PIXEL_SIZE && h_count < i_worm_x[3665:3660] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3665:3660] * PIXEL_SIZE && v_count < i_worm_y[3665:3660] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (611 < i_size && h_count >= i_worm_x[3671:3666] * PIXEL_SIZE && h_count < i_worm_x[3671:3666] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3671:3666] * PIXEL_SIZE && v_count < i_worm_y[3671:3666] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (612 < i_size && h_count >= i_worm_x[3677:3672] * PIXEL_SIZE && h_count < i_worm_x[3677:3672] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3677:3672] * PIXEL_SIZE && v_count < i_worm_y[3677:3672] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (613 < i_size && h_count >= i_worm_x[3683:3678] * PIXEL_SIZE && h_count < i_worm_x[3683:3678] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3683:3678] * PIXEL_SIZE && v_count < i_worm_y[3683:3678] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (614 < i_size && h_count >= i_worm_x[3689:3684] * PIXEL_SIZE && h_count < i_worm_x[3689:3684] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3689:3684] * PIXEL_SIZE && v_count < i_worm_y[3689:3684] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (615 < i_size && h_count >= i_worm_x[3695:3690] * PIXEL_SIZE && h_count < i_worm_x[3695:3690] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3695:3690] * PIXEL_SIZE && v_count < i_worm_y[3695:3690] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (616 < i_size && h_count >= i_worm_x[3701:3696] * PIXEL_SIZE && h_count < i_worm_x[3701:3696] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3701:3696] * PIXEL_SIZE && v_count < i_worm_y[3701:3696] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (617 < i_size && h_count >= i_worm_x[3707:3702] * PIXEL_SIZE && h_count < i_worm_x[3707:3702] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3707:3702] * PIXEL_SIZE && v_count < i_worm_y[3707:3702] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (618 < i_size && h_count >= i_worm_x[3713:3708] * PIXEL_SIZE && h_count < i_worm_x[3713:3708] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3713:3708] * PIXEL_SIZE && v_count < i_worm_y[3713:3708] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (619 < i_size && h_count >= i_worm_x[3719:3714] * PIXEL_SIZE && h_count < i_worm_x[3719:3714] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3719:3714] * PIXEL_SIZE && v_count < i_worm_y[3719:3714] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (620 < i_size && h_count >= i_worm_x[3725:3720] * PIXEL_SIZE && h_count < i_worm_x[3725:3720] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3725:3720] * PIXEL_SIZE && v_count < i_worm_y[3725:3720] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (621 < i_size && h_count >= i_worm_x[3731:3726] * PIXEL_SIZE && h_count < i_worm_x[3731:3726] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3731:3726] * PIXEL_SIZE && v_count < i_worm_y[3731:3726] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (622 < i_size && h_count >= i_worm_x[3737:3732] * PIXEL_SIZE && h_count < i_worm_x[3737:3732] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3737:3732] * PIXEL_SIZE && v_count < i_worm_y[3737:3732] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (623 < i_size && h_count >= i_worm_x[3743:3738] * PIXEL_SIZE && h_count < i_worm_x[3743:3738] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3743:3738] * PIXEL_SIZE && v_count < i_worm_y[3743:3738] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (624 < i_size && h_count >= i_worm_x[3749:3744] * PIXEL_SIZE && h_count < i_worm_x[3749:3744] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3749:3744] * PIXEL_SIZE && v_count < i_worm_y[3749:3744] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (625 < i_size && h_count >= i_worm_x[3755:3750] * PIXEL_SIZE && h_count < i_worm_x[3755:3750] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3755:3750] * PIXEL_SIZE && v_count < i_worm_y[3755:3750] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (626 < i_size && h_count >= i_worm_x[3761:3756] * PIXEL_SIZE && h_count < i_worm_x[3761:3756] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3761:3756] * PIXEL_SIZE && v_count < i_worm_y[3761:3756] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (627 < i_size && h_count >= i_worm_x[3767:3762] * PIXEL_SIZE && h_count < i_worm_x[3767:3762] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3767:3762] * PIXEL_SIZE && v_count < i_worm_y[3767:3762] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (628 < i_size && h_count >= i_worm_x[3773:3768] * PIXEL_SIZE && h_count < i_worm_x[3773:3768] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3773:3768] * PIXEL_SIZE && v_count < i_worm_y[3773:3768] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (629 < i_size && h_count >= i_worm_x[3779:3774] * PIXEL_SIZE && h_count < i_worm_x[3779:3774] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3779:3774] * PIXEL_SIZE && v_count < i_worm_y[3779:3774] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (630 < i_size && h_count >= i_worm_x[3785:3780] * PIXEL_SIZE && h_count < i_worm_x[3785:3780] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3785:3780] * PIXEL_SIZE && v_count < i_worm_y[3785:3780] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (631 < i_size && h_count >= i_worm_x[3791:3786] * PIXEL_SIZE && h_count < i_worm_x[3791:3786] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3791:3786] * PIXEL_SIZE && v_count < i_worm_y[3791:3786] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (632 < i_size && h_count >= i_worm_x[3797:3792] * PIXEL_SIZE && h_count < i_worm_x[3797:3792] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3797:3792] * PIXEL_SIZE && v_count < i_worm_y[3797:3792] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (633 < i_size && h_count >= i_worm_x[3803:3798] * PIXEL_SIZE && h_count < i_worm_x[3803:3798] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3803:3798] * PIXEL_SIZE && v_count < i_worm_y[3803:3798] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (634 < i_size && h_count >= i_worm_x[3809:3804] * PIXEL_SIZE && h_count < i_worm_x[3809:3804] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3809:3804] * PIXEL_SIZE && v_count < i_worm_y[3809:3804] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (635 < i_size && h_count >= i_worm_x[3815:3810] * PIXEL_SIZE && h_count < i_worm_x[3815:3810] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3815:3810] * PIXEL_SIZE && v_count < i_worm_y[3815:3810] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (636 < i_size && h_count >= i_worm_x[3821:3816] * PIXEL_SIZE && h_count < i_worm_x[3821:3816] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3821:3816] * PIXEL_SIZE && v_count < i_worm_y[3821:3816] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (637 < i_size && h_count >= i_worm_x[3827:3822] * PIXEL_SIZE && h_count < i_worm_x[3827:3822] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3827:3822] * PIXEL_SIZE && v_count < i_worm_y[3827:3822] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (638 < i_size && h_count >= i_worm_x[3833:3828] * PIXEL_SIZE && h_count < i_worm_x[3833:3828] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3833:3828] * PIXEL_SIZE && v_count < i_worm_y[3833:3828] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (639 < i_size && h_count >= i_worm_x[3839:3834] * PIXEL_SIZE && h_count < i_worm_x[3839:3834] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3839:3834] * PIXEL_SIZE && v_count < i_worm_y[3839:3834] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (640 < i_size && h_count >= i_worm_x[3845:3840] * PIXEL_SIZE && h_count < i_worm_x[3845:3840] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3845:3840] * PIXEL_SIZE && v_count < i_worm_y[3845:3840] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (641 < i_size && h_count >= i_worm_x[3851:3846] * PIXEL_SIZE && h_count < i_worm_x[3851:3846] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3851:3846] * PIXEL_SIZE && v_count < i_worm_y[3851:3846] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (642 < i_size && h_count >= i_worm_x[3857:3852] * PIXEL_SIZE && h_count < i_worm_x[3857:3852] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3857:3852] * PIXEL_SIZE && v_count < i_worm_y[3857:3852] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (643 < i_size && h_count >= i_worm_x[3863:3858] * PIXEL_SIZE && h_count < i_worm_x[3863:3858] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3863:3858] * PIXEL_SIZE && v_count < i_worm_y[3863:3858] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (644 < i_size && h_count >= i_worm_x[3869:3864] * PIXEL_SIZE && h_count < i_worm_x[3869:3864] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3869:3864] * PIXEL_SIZE && v_count < i_worm_y[3869:3864] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (645 < i_size && h_count >= i_worm_x[3875:3870] * PIXEL_SIZE && h_count < i_worm_x[3875:3870] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3875:3870] * PIXEL_SIZE && v_count < i_worm_y[3875:3870] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (646 < i_size && h_count >= i_worm_x[3881:3876] * PIXEL_SIZE && h_count < i_worm_x[3881:3876] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3881:3876] * PIXEL_SIZE && v_count < i_worm_y[3881:3876] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (647 < i_size && h_count >= i_worm_x[3887:3882] * PIXEL_SIZE && h_count < i_worm_x[3887:3882] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3887:3882] * PIXEL_SIZE && v_count < i_worm_y[3887:3882] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (648 < i_size && h_count >= i_worm_x[3893:3888] * PIXEL_SIZE && h_count < i_worm_x[3893:3888] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3893:3888] * PIXEL_SIZE && v_count < i_worm_y[3893:3888] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (649 < i_size && h_count >= i_worm_x[3899:3894] * PIXEL_SIZE && h_count < i_worm_x[3899:3894] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3899:3894] * PIXEL_SIZE && v_count < i_worm_y[3899:3894] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (650 < i_size && h_count >= i_worm_x[3905:3900] * PIXEL_SIZE && h_count < i_worm_x[3905:3900] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3905:3900] * PIXEL_SIZE && v_count < i_worm_y[3905:3900] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (651 < i_size && h_count >= i_worm_x[3911:3906] * PIXEL_SIZE && h_count < i_worm_x[3911:3906] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3911:3906] * PIXEL_SIZE && v_count < i_worm_y[3911:3906] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (652 < i_size && h_count >= i_worm_x[3917:3912] * PIXEL_SIZE && h_count < i_worm_x[3917:3912] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3917:3912] * PIXEL_SIZE && v_count < i_worm_y[3917:3912] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (653 < i_size && h_count >= i_worm_x[3923:3918] * PIXEL_SIZE && h_count < i_worm_x[3923:3918] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3923:3918] * PIXEL_SIZE && v_count < i_worm_y[3923:3918] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (654 < i_size && h_count >= i_worm_x[3929:3924] * PIXEL_SIZE && h_count < i_worm_x[3929:3924] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3929:3924] * PIXEL_SIZE && v_count < i_worm_y[3929:3924] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (655 < i_size && h_count >= i_worm_x[3935:3930] * PIXEL_SIZE && h_count < i_worm_x[3935:3930] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3935:3930] * PIXEL_SIZE && v_count < i_worm_y[3935:3930] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (656 < i_size && h_count >= i_worm_x[3941:3936] * PIXEL_SIZE && h_count < i_worm_x[3941:3936] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3941:3936] * PIXEL_SIZE && v_count < i_worm_y[3941:3936] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (657 < i_size && h_count >= i_worm_x[3947:3942] * PIXEL_SIZE && h_count < i_worm_x[3947:3942] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3947:3942] * PIXEL_SIZE && v_count < i_worm_y[3947:3942] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (658 < i_size && h_count >= i_worm_x[3953:3948] * PIXEL_SIZE && h_count < i_worm_x[3953:3948] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3953:3948] * PIXEL_SIZE && v_count < i_worm_y[3953:3948] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (659 < i_size && h_count >= i_worm_x[3959:3954] * PIXEL_SIZE && h_count < i_worm_x[3959:3954] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3959:3954] * PIXEL_SIZE && v_count < i_worm_y[3959:3954] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (660 < i_size && h_count >= i_worm_x[3965:3960] * PIXEL_SIZE && h_count < i_worm_x[3965:3960] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3965:3960] * PIXEL_SIZE && v_count < i_worm_y[3965:3960] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (661 < i_size && h_count >= i_worm_x[3971:3966] * PIXEL_SIZE && h_count < i_worm_x[3971:3966] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3971:3966] * PIXEL_SIZE && v_count < i_worm_y[3971:3966] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (662 < i_size && h_count >= i_worm_x[3977:3972] * PIXEL_SIZE && h_count < i_worm_x[3977:3972] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3977:3972] * PIXEL_SIZE && v_count < i_worm_y[3977:3972] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (663 < i_size && h_count >= i_worm_x[3983:3978] * PIXEL_SIZE && h_count < i_worm_x[3983:3978] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3983:3978] * PIXEL_SIZE && v_count < i_worm_y[3983:3978] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (664 < i_size && h_count >= i_worm_x[3989:3984] * PIXEL_SIZE && h_count < i_worm_x[3989:3984] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3989:3984] * PIXEL_SIZE && v_count < i_worm_y[3989:3984] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (665 < i_size && h_count >= i_worm_x[3995:3990] * PIXEL_SIZE && h_count < i_worm_x[3995:3990] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[3995:3990] * PIXEL_SIZE && v_count < i_worm_y[3995:3990] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (666 < i_size && h_count >= i_worm_x[4001:3996] * PIXEL_SIZE && h_count < i_worm_x[4001:3996] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4001:3996] * PIXEL_SIZE && v_count < i_worm_y[4001:3996] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (667 < i_size && h_count >= i_worm_x[4007:4002] * PIXEL_SIZE && h_count < i_worm_x[4007:4002] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4007:4002] * PIXEL_SIZE && v_count < i_worm_y[4007:4002] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (668 < i_size && h_count >= i_worm_x[4013:4008] * PIXEL_SIZE && h_count < i_worm_x[4013:4008] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4013:4008] * PIXEL_SIZE && v_count < i_worm_y[4013:4008] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (669 < i_size && h_count >= i_worm_x[4019:4014] * PIXEL_SIZE && h_count < i_worm_x[4019:4014] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4019:4014] * PIXEL_SIZE && v_count < i_worm_y[4019:4014] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (670 < i_size && h_count >= i_worm_x[4025:4020] * PIXEL_SIZE && h_count < i_worm_x[4025:4020] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4025:4020] * PIXEL_SIZE && v_count < i_worm_y[4025:4020] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (671 < i_size && h_count >= i_worm_x[4031:4026] * PIXEL_SIZE && h_count < i_worm_x[4031:4026] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4031:4026] * PIXEL_SIZE && v_count < i_worm_y[4031:4026] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (672 < i_size && h_count >= i_worm_x[4037:4032] * PIXEL_SIZE && h_count < i_worm_x[4037:4032] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4037:4032] * PIXEL_SIZE && v_count < i_worm_y[4037:4032] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (673 < i_size && h_count >= i_worm_x[4043:4038] * PIXEL_SIZE && h_count < i_worm_x[4043:4038] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4043:4038] * PIXEL_SIZE && v_count < i_worm_y[4043:4038] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (674 < i_size && h_count >= i_worm_x[4049:4044] * PIXEL_SIZE && h_count < i_worm_x[4049:4044] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4049:4044] * PIXEL_SIZE && v_count < i_worm_y[4049:4044] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (675 < i_size && h_count >= i_worm_x[4055:4050] * PIXEL_SIZE && h_count < i_worm_x[4055:4050] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4055:4050] * PIXEL_SIZE && v_count < i_worm_y[4055:4050] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (676 < i_size && h_count >= i_worm_x[4061:4056] * PIXEL_SIZE && h_count < i_worm_x[4061:4056] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4061:4056] * PIXEL_SIZE && v_count < i_worm_y[4061:4056] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (677 < i_size && h_count >= i_worm_x[4067:4062] * PIXEL_SIZE && h_count < i_worm_x[4067:4062] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4067:4062] * PIXEL_SIZE && v_count < i_worm_y[4067:4062] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (678 < i_size && h_count >= i_worm_x[4073:4068] * PIXEL_SIZE && h_count < i_worm_x[4073:4068] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4073:4068] * PIXEL_SIZE && v_count < i_worm_y[4073:4068] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (679 < i_size && h_count >= i_worm_x[4079:4074] * PIXEL_SIZE && h_count < i_worm_x[4079:4074] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4079:4074] * PIXEL_SIZE && v_count < i_worm_y[4079:4074] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (680 < i_size && h_count >= i_worm_x[4085:4080] * PIXEL_SIZE && h_count < i_worm_x[4085:4080] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4085:4080] * PIXEL_SIZE && v_count < i_worm_y[4085:4080] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (681 < i_size && h_count >= i_worm_x[4091:4086] * PIXEL_SIZE && h_count < i_worm_x[4091:4086] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4091:4086] * PIXEL_SIZE && v_count < i_worm_y[4091:4086] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (682 < i_size && h_count >= i_worm_x[4097:4092] * PIXEL_SIZE && h_count < i_worm_x[4097:4092] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4097:4092] * PIXEL_SIZE && v_count < i_worm_y[4097:4092] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (683 < i_size && h_count >= i_worm_x[4103:4098] * PIXEL_SIZE && h_count < i_worm_x[4103:4098] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4103:4098] * PIXEL_SIZE && v_count < i_worm_y[4103:4098] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (684 < i_size && h_count >= i_worm_x[4109:4104] * PIXEL_SIZE && h_count < i_worm_x[4109:4104] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4109:4104] * PIXEL_SIZE && v_count < i_worm_y[4109:4104] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (685 < i_size && h_count >= i_worm_x[4115:4110] * PIXEL_SIZE && h_count < i_worm_x[4115:4110] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4115:4110] * PIXEL_SIZE && v_count < i_worm_y[4115:4110] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (686 < i_size && h_count >= i_worm_x[4121:4116] * PIXEL_SIZE && h_count < i_worm_x[4121:4116] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4121:4116] * PIXEL_SIZE && v_count < i_worm_y[4121:4116] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (687 < i_size && h_count >= i_worm_x[4127:4122] * PIXEL_SIZE && h_count < i_worm_x[4127:4122] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4127:4122] * PIXEL_SIZE && v_count < i_worm_y[4127:4122] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (688 < i_size && h_count >= i_worm_x[4133:4128] * PIXEL_SIZE && h_count < i_worm_x[4133:4128] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4133:4128] * PIXEL_SIZE && v_count < i_worm_y[4133:4128] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (689 < i_size && h_count >= i_worm_x[4139:4134] * PIXEL_SIZE && h_count < i_worm_x[4139:4134] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4139:4134] * PIXEL_SIZE && v_count < i_worm_y[4139:4134] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (690 < i_size && h_count >= i_worm_x[4145:4140] * PIXEL_SIZE && h_count < i_worm_x[4145:4140] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4145:4140] * PIXEL_SIZE && v_count < i_worm_y[4145:4140] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (691 < i_size && h_count >= i_worm_x[4151:4146] * PIXEL_SIZE && h_count < i_worm_x[4151:4146] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4151:4146] * PIXEL_SIZE && v_count < i_worm_y[4151:4146] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (692 < i_size && h_count >= i_worm_x[4157:4152] * PIXEL_SIZE && h_count < i_worm_x[4157:4152] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4157:4152] * PIXEL_SIZE && v_count < i_worm_y[4157:4152] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (693 < i_size && h_count >= i_worm_x[4163:4158] * PIXEL_SIZE && h_count < i_worm_x[4163:4158] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4163:4158] * PIXEL_SIZE && v_count < i_worm_y[4163:4158] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (694 < i_size && h_count >= i_worm_x[4169:4164] * PIXEL_SIZE && h_count < i_worm_x[4169:4164] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4169:4164] * PIXEL_SIZE && v_count < i_worm_y[4169:4164] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (695 < i_size && h_count >= i_worm_x[4175:4170] * PIXEL_SIZE && h_count < i_worm_x[4175:4170] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4175:4170] * PIXEL_SIZE && v_count < i_worm_y[4175:4170] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (696 < i_size && h_count >= i_worm_x[4181:4176] * PIXEL_SIZE && h_count < i_worm_x[4181:4176] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4181:4176] * PIXEL_SIZE && v_count < i_worm_y[4181:4176] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (697 < i_size && h_count >= i_worm_x[4187:4182] * PIXEL_SIZE && h_count < i_worm_x[4187:4182] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4187:4182] * PIXEL_SIZE && v_count < i_worm_y[4187:4182] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (698 < i_size && h_count >= i_worm_x[4193:4188] * PIXEL_SIZE && h_count < i_worm_x[4193:4188] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4193:4188] * PIXEL_SIZE && v_count < i_worm_y[4193:4188] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (699 < i_size && h_count >= i_worm_x[4199:4194] * PIXEL_SIZE && h_count < i_worm_x[4199:4194] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4199:4194] * PIXEL_SIZE && v_count < i_worm_y[4199:4194] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (700 < i_size && h_count >= i_worm_x[4205:4200] * PIXEL_SIZE && h_count < i_worm_x[4205:4200] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4205:4200] * PIXEL_SIZE && v_count < i_worm_y[4205:4200] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (701 < i_size && h_count >= i_worm_x[4211:4206] * PIXEL_SIZE && h_count < i_worm_x[4211:4206] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4211:4206] * PIXEL_SIZE && v_count < i_worm_y[4211:4206] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (702 < i_size && h_count >= i_worm_x[4217:4212] * PIXEL_SIZE && h_count < i_worm_x[4217:4212] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4217:4212] * PIXEL_SIZE && v_count < i_worm_y[4217:4212] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (703 < i_size && h_count >= i_worm_x[4223:4218] * PIXEL_SIZE && h_count < i_worm_x[4223:4218] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4223:4218] * PIXEL_SIZE && v_count < i_worm_y[4223:4218] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (704 < i_size && h_count >= i_worm_x[4229:4224] * PIXEL_SIZE && h_count < i_worm_x[4229:4224] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4229:4224] * PIXEL_SIZE && v_count < i_worm_y[4229:4224] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (705 < i_size && h_count >= i_worm_x[4235:4230] * PIXEL_SIZE && h_count < i_worm_x[4235:4230] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4235:4230] * PIXEL_SIZE && v_count < i_worm_y[4235:4230] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (706 < i_size && h_count >= i_worm_x[4241:4236] * PIXEL_SIZE && h_count < i_worm_x[4241:4236] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4241:4236] * PIXEL_SIZE && v_count < i_worm_y[4241:4236] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (707 < i_size && h_count >= i_worm_x[4247:4242] * PIXEL_SIZE && h_count < i_worm_x[4247:4242] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4247:4242] * PIXEL_SIZE && v_count < i_worm_y[4247:4242] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (708 < i_size && h_count >= i_worm_x[4253:4248] * PIXEL_SIZE && h_count < i_worm_x[4253:4248] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4253:4248] * PIXEL_SIZE && v_count < i_worm_y[4253:4248] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (709 < i_size && h_count >= i_worm_x[4259:4254] * PIXEL_SIZE && h_count < i_worm_x[4259:4254] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4259:4254] * PIXEL_SIZE && v_count < i_worm_y[4259:4254] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (710 < i_size && h_count >= i_worm_x[4265:4260] * PIXEL_SIZE && h_count < i_worm_x[4265:4260] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4265:4260] * PIXEL_SIZE && v_count < i_worm_y[4265:4260] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (711 < i_size && h_count >= i_worm_x[4271:4266] * PIXEL_SIZE && h_count < i_worm_x[4271:4266] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4271:4266] * PIXEL_SIZE && v_count < i_worm_y[4271:4266] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (712 < i_size && h_count >= i_worm_x[4277:4272] * PIXEL_SIZE && h_count < i_worm_x[4277:4272] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4277:4272] * PIXEL_SIZE && v_count < i_worm_y[4277:4272] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (713 < i_size && h_count >= i_worm_x[4283:4278] * PIXEL_SIZE && h_count < i_worm_x[4283:4278] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4283:4278] * PIXEL_SIZE && v_count < i_worm_y[4283:4278] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (714 < i_size && h_count >= i_worm_x[4289:4284] * PIXEL_SIZE && h_count < i_worm_x[4289:4284] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4289:4284] * PIXEL_SIZE && v_count < i_worm_y[4289:4284] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (715 < i_size && h_count >= i_worm_x[4295:4290] * PIXEL_SIZE && h_count < i_worm_x[4295:4290] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4295:4290] * PIXEL_SIZE && v_count < i_worm_y[4295:4290] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (716 < i_size && h_count >= i_worm_x[4301:4296] * PIXEL_SIZE && h_count < i_worm_x[4301:4296] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4301:4296] * PIXEL_SIZE && v_count < i_worm_y[4301:4296] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (717 < i_size && h_count >= i_worm_x[4307:4302] * PIXEL_SIZE && h_count < i_worm_x[4307:4302] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4307:4302] * PIXEL_SIZE && v_count < i_worm_y[4307:4302] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (718 < i_size && h_count >= i_worm_x[4313:4308] * PIXEL_SIZE && h_count < i_worm_x[4313:4308] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4313:4308] * PIXEL_SIZE && v_count < i_worm_y[4313:4308] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (719 < i_size && h_count >= i_worm_x[4319:4314] * PIXEL_SIZE && h_count < i_worm_x[4319:4314] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4319:4314] * PIXEL_SIZE && v_count < i_worm_y[4319:4314] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (720 < i_size && h_count >= i_worm_x[4325:4320] * PIXEL_SIZE && h_count < i_worm_x[4325:4320] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4325:4320] * PIXEL_SIZE && v_count < i_worm_y[4325:4320] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (721 < i_size && h_count >= i_worm_x[4331:4326] * PIXEL_SIZE && h_count < i_worm_x[4331:4326] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4331:4326] * PIXEL_SIZE && v_count < i_worm_y[4331:4326] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (722 < i_size && h_count >= i_worm_x[4337:4332] * PIXEL_SIZE && h_count < i_worm_x[4337:4332] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4337:4332] * PIXEL_SIZE && v_count < i_worm_y[4337:4332] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (723 < i_size && h_count >= i_worm_x[4343:4338] * PIXEL_SIZE && h_count < i_worm_x[4343:4338] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4343:4338] * PIXEL_SIZE && v_count < i_worm_y[4343:4338] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (724 < i_size && h_count >= i_worm_x[4349:4344] * PIXEL_SIZE && h_count < i_worm_x[4349:4344] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4349:4344] * PIXEL_SIZE && v_count < i_worm_y[4349:4344] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (725 < i_size && h_count >= i_worm_x[4355:4350] * PIXEL_SIZE && h_count < i_worm_x[4355:4350] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4355:4350] * PIXEL_SIZE && v_count < i_worm_y[4355:4350] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (726 < i_size && h_count >= i_worm_x[4361:4356] * PIXEL_SIZE && h_count < i_worm_x[4361:4356] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4361:4356] * PIXEL_SIZE && v_count < i_worm_y[4361:4356] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (727 < i_size && h_count >= i_worm_x[4367:4362] * PIXEL_SIZE && h_count < i_worm_x[4367:4362] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4367:4362] * PIXEL_SIZE && v_count < i_worm_y[4367:4362] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (728 < i_size && h_count >= i_worm_x[4373:4368] * PIXEL_SIZE && h_count < i_worm_x[4373:4368] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4373:4368] * PIXEL_SIZE && v_count < i_worm_y[4373:4368] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (729 < i_size && h_count >= i_worm_x[4379:4374] * PIXEL_SIZE && h_count < i_worm_x[4379:4374] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4379:4374] * PIXEL_SIZE && v_count < i_worm_y[4379:4374] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (730 < i_size && h_count >= i_worm_x[4385:4380] * PIXEL_SIZE && h_count < i_worm_x[4385:4380] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4385:4380] * PIXEL_SIZE && v_count < i_worm_y[4385:4380] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (731 < i_size && h_count >= i_worm_x[4391:4386] * PIXEL_SIZE && h_count < i_worm_x[4391:4386] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4391:4386] * PIXEL_SIZE && v_count < i_worm_y[4391:4386] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (732 < i_size && h_count >= i_worm_x[4397:4392] * PIXEL_SIZE && h_count < i_worm_x[4397:4392] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4397:4392] * PIXEL_SIZE && v_count < i_worm_y[4397:4392] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (733 < i_size && h_count >= i_worm_x[4403:4398] * PIXEL_SIZE && h_count < i_worm_x[4403:4398] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4403:4398] * PIXEL_SIZE && v_count < i_worm_y[4403:4398] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (734 < i_size && h_count >= i_worm_x[4409:4404] * PIXEL_SIZE && h_count < i_worm_x[4409:4404] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4409:4404] * PIXEL_SIZE && v_count < i_worm_y[4409:4404] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (735 < i_size && h_count >= i_worm_x[4415:4410] * PIXEL_SIZE && h_count < i_worm_x[4415:4410] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4415:4410] * PIXEL_SIZE && v_count < i_worm_y[4415:4410] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (736 < i_size && h_count >= i_worm_x[4421:4416] * PIXEL_SIZE && h_count < i_worm_x[4421:4416] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4421:4416] * PIXEL_SIZE && v_count < i_worm_y[4421:4416] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (737 < i_size && h_count >= i_worm_x[4427:4422] * PIXEL_SIZE && h_count < i_worm_x[4427:4422] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4427:4422] * PIXEL_SIZE && v_count < i_worm_y[4427:4422] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (738 < i_size && h_count >= i_worm_x[4433:4428] * PIXEL_SIZE && h_count < i_worm_x[4433:4428] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4433:4428] * PIXEL_SIZE && v_count < i_worm_y[4433:4428] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (739 < i_size && h_count >= i_worm_x[4439:4434] * PIXEL_SIZE && h_count < i_worm_x[4439:4434] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4439:4434] * PIXEL_SIZE && v_count < i_worm_y[4439:4434] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (740 < i_size && h_count >= i_worm_x[4445:4440] * PIXEL_SIZE && h_count < i_worm_x[4445:4440] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4445:4440] * PIXEL_SIZE && v_count < i_worm_y[4445:4440] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (741 < i_size && h_count >= i_worm_x[4451:4446] * PIXEL_SIZE && h_count < i_worm_x[4451:4446] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4451:4446] * PIXEL_SIZE && v_count < i_worm_y[4451:4446] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (742 < i_size && h_count >= i_worm_x[4457:4452] * PIXEL_SIZE && h_count < i_worm_x[4457:4452] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4457:4452] * PIXEL_SIZE && v_count < i_worm_y[4457:4452] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (743 < i_size && h_count >= i_worm_x[4463:4458] * PIXEL_SIZE && h_count < i_worm_x[4463:4458] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4463:4458] * PIXEL_SIZE && v_count < i_worm_y[4463:4458] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (744 < i_size && h_count >= i_worm_x[4469:4464] * PIXEL_SIZE && h_count < i_worm_x[4469:4464] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4469:4464] * PIXEL_SIZE && v_count < i_worm_y[4469:4464] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (745 < i_size && h_count >= i_worm_x[4475:4470] * PIXEL_SIZE && h_count < i_worm_x[4475:4470] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4475:4470] * PIXEL_SIZE && v_count < i_worm_y[4475:4470] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (746 < i_size && h_count >= i_worm_x[4481:4476] * PIXEL_SIZE && h_count < i_worm_x[4481:4476] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4481:4476] * PIXEL_SIZE && v_count < i_worm_y[4481:4476] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (747 < i_size && h_count >= i_worm_x[4487:4482] * PIXEL_SIZE && h_count < i_worm_x[4487:4482] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4487:4482] * PIXEL_SIZE && v_count < i_worm_y[4487:4482] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (748 < i_size && h_count >= i_worm_x[4493:4488] * PIXEL_SIZE && h_count < i_worm_x[4493:4488] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4493:4488] * PIXEL_SIZE && v_count < i_worm_y[4493:4488] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (749 < i_size && h_count >= i_worm_x[4499:4494] * PIXEL_SIZE && h_count < i_worm_x[4499:4494] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4499:4494] * PIXEL_SIZE && v_count < i_worm_y[4499:4494] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (750 < i_size && h_count >= i_worm_x[4505:4500] * PIXEL_SIZE && h_count < i_worm_x[4505:4500] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4505:4500] * PIXEL_SIZE && v_count < i_worm_y[4505:4500] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (751 < i_size && h_count >= i_worm_x[4511:4506] * PIXEL_SIZE && h_count < i_worm_x[4511:4506] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4511:4506] * PIXEL_SIZE && v_count < i_worm_y[4511:4506] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (752 < i_size && h_count >= i_worm_x[4517:4512] * PIXEL_SIZE && h_count < i_worm_x[4517:4512] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4517:4512] * PIXEL_SIZE && v_count < i_worm_y[4517:4512] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (753 < i_size && h_count >= i_worm_x[4523:4518] * PIXEL_SIZE && h_count < i_worm_x[4523:4518] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4523:4518] * PIXEL_SIZE && v_count < i_worm_y[4523:4518] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (754 < i_size && h_count >= i_worm_x[4529:4524] * PIXEL_SIZE && h_count < i_worm_x[4529:4524] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4529:4524] * PIXEL_SIZE && v_count < i_worm_y[4529:4524] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (755 < i_size && h_count >= i_worm_x[4535:4530] * PIXEL_SIZE && h_count < i_worm_x[4535:4530] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4535:4530] * PIXEL_SIZE && v_count < i_worm_y[4535:4530] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (756 < i_size && h_count >= i_worm_x[4541:4536] * PIXEL_SIZE && h_count < i_worm_x[4541:4536] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4541:4536] * PIXEL_SIZE && v_count < i_worm_y[4541:4536] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (757 < i_size && h_count >= i_worm_x[4547:4542] * PIXEL_SIZE && h_count < i_worm_x[4547:4542] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4547:4542] * PIXEL_SIZE && v_count < i_worm_y[4547:4542] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (758 < i_size && h_count >= i_worm_x[4553:4548] * PIXEL_SIZE && h_count < i_worm_x[4553:4548] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4553:4548] * PIXEL_SIZE && v_count < i_worm_y[4553:4548] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (759 < i_size && h_count >= i_worm_x[4559:4554] * PIXEL_SIZE && h_count < i_worm_x[4559:4554] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4559:4554] * PIXEL_SIZE && v_count < i_worm_y[4559:4554] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (760 < i_size && h_count >= i_worm_x[4565:4560] * PIXEL_SIZE && h_count < i_worm_x[4565:4560] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4565:4560] * PIXEL_SIZE && v_count < i_worm_y[4565:4560] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (761 < i_size && h_count >= i_worm_x[4571:4566] * PIXEL_SIZE && h_count < i_worm_x[4571:4566] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4571:4566] * PIXEL_SIZE && v_count < i_worm_y[4571:4566] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (762 < i_size && h_count >= i_worm_x[4577:4572] * PIXEL_SIZE && h_count < i_worm_x[4577:4572] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4577:4572] * PIXEL_SIZE && v_count < i_worm_y[4577:4572] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (763 < i_size && h_count >= i_worm_x[4583:4578] * PIXEL_SIZE && h_count < i_worm_x[4583:4578] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4583:4578] * PIXEL_SIZE && v_count < i_worm_y[4583:4578] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (764 < i_size && h_count >= i_worm_x[4589:4584] * PIXEL_SIZE && h_count < i_worm_x[4589:4584] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4589:4584] * PIXEL_SIZE && v_count < i_worm_y[4589:4584] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (765 < i_size && h_count >= i_worm_x[4595:4590] * PIXEL_SIZE && h_count < i_worm_x[4595:4590] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4595:4590] * PIXEL_SIZE && v_count < i_worm_y[4595:4590] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (766 < i_size && h_count >= i_worm_x[4601:4596] * PIXEL_SIZE && h_count < i_worm_x[4601:4596] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4601:4596] * PIXEL_SIZE && v_count < i_worm_y[4601:4596] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (767 < i_size && h_count >= i_worm_x[4607:4602] * PIXEL_SIZE && h_count < i_worm_x[4607:4602] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4607:4602] * PIXEL_SIZE && v_count < i_worm_y[4607:4602] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (768 < i_size && h_count >= i_worm_x[4613:4608] * PIXEL_SIZE && h_count < i_worm_x[4613:4608] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4613:4608] * PIXEL_SIZE && v_count < i_worm_y[4613:4608] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (769 < i_size && h_count >= i_worm_x[4619:4614] * PIXEL_SIZE && h_count < i_worm_x[4619:4614] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4619:4614] * PIXEL_SIZE && v_count < i_worm_y[4619:4614] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (770 < i_size && h_count >= i_worm_x[4625:4620] * PIXEL_SIZE && h_count < i_worm_x[4625:4620] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4625:4620] * PIXEL_SIZE && v_count < i_worm_y[4625:4620] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (771 < i_size && h_count >= i_worm_x[4631:4626] * PIXEL_SIZE && h_count < i_worm_x[4631:4626] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4631:4626] * PIXEL_SIZE && v_count < i_worm_y[4631:4626] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (772 < i_size && h_count >= i_worm_x[4637:4632] * PIXEL_SIZE && h_count < i_worm_x[4637:4632] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4637:4632] * PIXEL_SIZE && v_count < i_worm_y[4637:4632] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (773 < i_size && h_count >= i_worm_x[4643:4638] * PIXEL_SIZE && h_count < i_worm_x[4643:4638] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4643:4638] * PIXEL_SIZE && v_count < i_worm_y[4643:4638] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (774 < i_size && h_count >= i_worm_x[4649:4644] * PIXEL_SIZE && h_count < i_worm_x[4649:4644] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4649:4644] * PIXEL_SIZE && v_count < i_worm_y[4649:4644] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (775 < i_size && h_count >= i_worm_x[4655:4650] * PIXEL_SIZE && h_count < i_worm_x[4655:4650] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4655:4650] * PIXEL_SIZE && v_count < i_worm_y[4655:4650] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (776 < i_size && h_count >= i_worm_x[4661:4656] * PIXEL_SIZE && h_count < i_worm_x[4661:4656] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4661:4656] * PIXEL_SIZE && v_count < i_worm_y[4661:4656] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (777 < i_size && h_count >= i_worm_x[4667:4662] * PIXEL_SIZE && h_count < i_worm_x[4667:4662] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4667:4662] * PIXEL_SIZE && v_count < i_worm_y[4667:4662] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (778 < i_size && h_count >= i_worm_x[4673:4668] * PIXEL_SIZE && h_count < i_worm_x[4673:4668] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4673:4668] * PIXEL_SIZE && v_count < i_worm_y[4673:4668] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (779 < i_size && h_count >= i_worm_x[4679:4674] * PIXEL_SIZE && h_count < i_worm_x[4679:4674] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4679:4674] * PIXEL_SIZE && v_count < i_worm_y[4679:4674] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (780 < i_size && h_count >= i_worm_x[4685:4680] * PIXEL_SIZE && h_count < i_worm_x[4685:4680] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4685:4680] * PIXEL_SIZE && v_count < i_worm_y[4685:4680] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (781 < i_size && h_count >= i_worm_x[4691:4686] * PIXEL_SIZE && h_count < i_worm_x[4691:4686] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4691:4686] * PIXEL_SIZE && v_count < i_worm_y[4691:4686] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (782 < i_size && h_count >= i_worm_x[4697:4692] * PIXEL_SIZE && h_count < i_worm_x[4697:4692] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4697:4692] * PIXEL_SIZE && v_count < i_worm_y[4697:4692] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (783 < i_size && h_count >= i_worm_x[4703:4698] * PIXEL_SIZE && h_count < i_worm_x[4703:4698] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4703:4698] * PIXEL_SIZE && v_count < i_worm_y[4703:4698] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (784 < i_size && h_count >= i_worm_x[4709:4704] * PIXEL_SIZE && h_count < i_worm_x[4709:4704] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4709:4704] * PIXEL_SIZE && v_count < i_worm_y[4709:4704] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (785 < i_size && h_count >= i_worm_x[4715:4710] * PIXEL_SIZE && h_count < i_worm_x[4715:4710] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4715:4710] * PIXEL_SIZE && v_count < i_worm_y[4715:4710] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (786 < i_size && h_count >= i_worm_x[4721:4716] * PIXEL_SIZE && h_count < i_worm_x[4721:4716] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4721:4716] * PIXEL_SIZE && v_count < i_worm_y[4721:4716] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (787 < i_size && h_count >= i_worm_x[4727:4722] * PIXEL_SIZE && h_count < i_worm_x[4727:4722] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4727:4722] * PIXEL_SIZE && v_count < i_worm_y[4727:4722] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (788 < i_size && h_count >= i_worm_x[4733:4728] * PIXEL_SIZE && h_count < i_worm_x[4733:4728] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4733:4728] * PIXEL_SIZE && v_count < i_worm_y[4733:4728] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (789 < i_size && h_count >= i_worm_x[4739:4734] * PIXEL_SIZE && h_count < i_worm_x[4739:4734] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4739:4734] * PIXEL_SIZE && v_count < i_worm_y[4739:4734] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (790 < i_size && h_count >= i_worm_x[4745:4740] * PIXEL_SIZE && h_count < i_worm_x[4745:4740] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4745:4740] * PIXEL_SIZE && v_count < i_worm_y[4745:4740] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (791 < i_size && h_count >= i_worm_x[4751:4746] * PIXEL_SIZE && h_count < i_worm_x[4751:4746] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4751:4746] * PIXEL_SIZE && v_count < i_worm_y[4751:4746] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (792 < i_size && h_count >= i_worm_x[4757:4752] * PIXEL_SIZE && h_count < i_worm_x[4757:4752] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4757:4752] * PIXEL_SIZE && v_count < i_worm_y[4757:4752] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (793 < i_size && h_count >= i_worm_x[4763:4758] * PIXEL_SIZE && h_count < i_worm_x[4763:4758] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4763:4758] * PIXEL_SIZE && v_count < i_worm_y[4763:4758] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (794 < i_size && h_count >= i_worm_x[4769:4764] * PIXEL_SIZE && h_count < i_worm_x[4769:4764] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4769:4764] * PIXEL_SIZE && v_count < i_worm_y[4769:4764] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (795 < i_size && h_count >= i_worm_x[4775:4770] * PIXEL_SIZE && h_count < i_worm_x[4775:4770] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4775:4770] * PIXEL_SIZE && v_count < i_worm_y[4775:4770] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (796 < i_size && h_count >= i_worm_x[4781:4776] * PIXEL_SIZE && h_count < i_worm_x[4781:4776] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4781:4776] * PIXEL_SIZE && v_count < i_worm_y[4781:4776] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (797 < i_size && h_count >= i_worm_x[4787:4782] * PIXEL_SIZE && h_count < i_worm_x[4787:4782] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4787:4782] * PIXEL_SIZE && v_count < i_worm_y[4787:4782] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (798 < i_size && h_count >= i_worm_x[4793:4788] * PIXEL_SIZE && h_count < i_worm_x[4793:4788] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4793:4788] * PIXEL_SIZE && v_count < i_worm_y[4793:4788] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (799 < i_size && h_count >= i_worm_x[4799:4794] * PIXEL_SIZE && h_count < i_worm_x[4799:4794] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4799:4794] * PIXEL_SIZE && v_count < i_worm_y[4799:4794] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (800 < i_size && h_count >= i_worm_x[4805:4800] * PIXEL_SIZE && h_count < i_worm_x[4805:4800] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4805:4800] * PIXEL_SIZE && v_count < i_worm_y[4805:4800] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (801 < i_size && h_count >= i_worm_x[4811:4806] * PIXEL_SIZE && h_count < i_worm_x[4811:4806] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4811:4806] * PIXEL_SIZE && v_count < i_worm_y[4811:4806] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (802 < i_size && h_count >= i_worm_x[4817:4812] * PIXEL_SIZE && h_count < i_worm_x[4817:4812] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4817:4812] * PIXEL_SIZE && v_count < i_worm_y[4817:4812] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (803 < i_size && h_count >= i_worm_x[4823:4818] * PIXEL_SIZE && h_count < i_worm_x[4823:4818] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4823:4818] * PIXEL_SIZE && v_count < i_worm_y[4823:4818] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (804 < i_size && h_count >= i_worm_x[4829:4824] * PIXEL_SIZE && h_count < i_worm_x[4829:4824] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4829:4824] * PIXEL_SIZE && v_count < i_worm_y[4829:4824] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (805 < i_size && h_count >= i_worm_x[4835:4830] * PIXEL_SIZE && h_count < i_worm_x[4835:4830] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4835:4830] * PIXEL_SIZE && v_count < i_worm_y[4835:4830] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (806 < i_size && h_count >= i_worm_x[4841:4836] * PIXEL_SIZE && h_count < i_worm_x[4841:4836] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4841:4836] * PIXEL_SIZE && v_count < i_worm_y[4841:4836] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (807 < i_size && h_count >= i_worm_x[4847:4842] * PIXEL_SIZE && h_count < i_worm_x[4847:4842] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4847:4842] * PIXEL_SIZE && v_count < i_worm_y[4847:4842] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (808 < i_size && h_count >= i_worm_x[4853:4848] * PIXEL_SIZE && h_count < i_worm_x[4853:4848] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4853:4848] * PIXEL_SIZE && v_count < i_worm_y[4853:4848] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (809 < i_size && h_count >= i_worm_x[4859:4854] * PIXEL_SIZE && h_count < i_worm_x[4859:4854] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4859:4854] * PIXEL_SIZE && v_count < i_worm_y[4859:4854] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (810 < i_size && h_count >= i_worm_x[4865:4860] * PIXEL_SIZE && h_count < i_worm_x[4865:4860] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4865:4860] * PIXEL_SIZE && v_count < i_worm_y[4865:4860] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (811 < i_size && h_count >= i_worm_x[4871:4866] * PIXEL_SIZE && h_count < i_worm_x[4871:4866] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4871:4866] * PIXEL_SIZE && v_count < i_worm_y[4871:4866] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (812 < i_size && h_count >= i_worm_x[4877:4872] * PIXEL_SIZE && h_count < i_worm_x[4877:4872] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4877:4872] * PIXEL_SIZE && v_count < i_worm_y[4877:4872] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (813 < i_size && h_count >= i_worm_x[4883:4878] * PIXEL_SIZE && h_count < i_worm_x[4883:4878] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4883:4878] * PIXEL_SIZE && v_count < i_worm_y[4883:4878] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (814 < i_size && h_count >= i_worm_x[4889:4884] * PIXEL_SIZE && h_count < i_worm_x[4889:4884] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4889:4884] * PIXEL_SIZE && v_count < i_worm_y[4889:4884] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (815 < i_size && h_count >= i_worm_x[4895:4890] * PIXEL_SIZE && h_count < i_worm_x[4895:4890] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4895:4890] * PIXEL_SIZE && v_count < i_worm_y[4895:4890] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (816 < i_size && h_count >= i_worm_x[4901:4896] * PIXEL_SIZE && h_count < i_worm_x[4901:4896] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4901:4896] * PIXEL_SIZE && v_count < i_worm_y[4901:4896] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (817 < i_size && h_count >= i_worm_x[4907:4902] * PIXEL_SIZE && h_count < i_worm_x[4907:4902] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4907:4902] * PIXEL_SIZE && v_count < i_worm_y[4907:4902] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (818 < i_size && h_count >= i_worm_x[4913:4908] * PIXEL_SIZE && h_count < i_worm_x[4913:4908] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4913:4908] * PIXEL_SIZE && v_count < i_worm_y[4913:4908] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (819 < i_size && h_count >= i_worm_x[4919:4914] * PIXEL_SIZE && h_count < i_worm_x[4919:4914] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4919:4914] * PIXEL_SIZE && v_count < i_worm_y[4919:4914] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (820 < i_size && h_count >= i_worm_x[4925:4920] * PIXEL_SIZE && h_count < i_worm_x[4925:4920] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4925:4920] * PIXEL_SIZE && v_count < i_worm_y[4925:4920] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (821 < i_size && h_count >= i_worm_x[4931:4926] * PIXEL_SIZE && h_count < i_worm_x[4931:4926] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4931:4926] * PIXEL_SIZE && v_count < i_worm_y[4931:4926] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (822 < i_size && h_count >= i_worm_x[4937:4932] * PIXEL_SIZE && h_count < i_worm_x[4937:4932] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4937:4932] * PIXEL_SIZE && v_count < i_worm_y[4937:4932] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (823 < i_size && h_count >= i_worm_x[4943:4938] * PIXEL_SIZE && h_count < i_worm_x[4943:4938] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4943:4938] * PIXEL_SIZE && v_count < i_worm_y[4943:4938] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (824 < i_size && h_count >= i_worm_x[4949:4944] * PIXEL_SIZE && h_count < i_worm_x[4949:4944] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4949:4944] * PIXEL_SIZE && v_count < i_worm_y[4949:4944] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (825 < i_size && h_count >= i_worm_x[4955:4950] * PIXEL_SIZE && h_count < i_worm_x[4955:4950] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4955:4950] * PIXEL_SIZE && v_count < i_worm_y[4955:4950] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (826 < i_size && h_count >= i_worm_x[4961:4956] * PIXEL_SIZE && h_count < i_worm_x[4961:4956] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4961:4956] * PIXEL_SIZE && v_count < i_worm_y[4961:4956] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (827 < i_size && h_count >= i_worm_x[4967:4962] * PIXEL_SIZE && h_count < i_worm_x[4967:4962] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4967:4962] * PIXEL_SIZE && v_count < i_worm_y[4967:4962] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (828 < i_size && h_count >= i_worm_x[4973:4968] * PIXEL_SIZE && h_count < i_worm_x[4973:4968] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4973:4968] * PIXEL_SIZE && v_count < i_worm_y[4973:4968] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (829 < i_size && h_count >= i_worm_x[4979:4974] * PIXEL_SIZE && h_count < i_worm_x[4979:4974] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4979:4974] * PIXEL_SIZE && v_count < i_worm_y[4979:4974] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (830 < i_size && h_count >= i_worm_x[4985:4980] * PIXEL_SIZE && h_count < i_worm_x[4985:4980] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4985:4980] * PIXEL_SIZE && v_count < i_worm_y[4985:4980] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (831 < i_size && h_count >= i_worm_x[4991:4986] * PIXEL_SIZE && h_count < i_worm_x[4991:4986] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4991:4986] * PIXEL_SIZE && v_count < i_worm_y[4991:4986] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (832 < i_size && h_count >= i_worm_x[4997:4992] * PIXEL_SIZE && h_count < i_worm_x[4997:4992] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[4997:4992] * PIXEL_SIZE && v_count < i_worm_y[4997:4992] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (833 < i_size && h_count >= i_worm_x[5003:4998] * PIXEL_SIZE && h_count < i_worm_x[5003:4998] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5003:4998] * PIXEL_SIZE && v_count < i_worm_y[5003:4998] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (834 < i_size && h_count >= i_worm_x[5009:5004] * PIXEL_SIZE && h_count < i_worm_x[5009:5004] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5009:5004] * PIXEL_SIZE && v_count < i_worm_y[5009:5004] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (835 < i_size && h_count >= i_worm_x[5015:5010] * PIXEL_SIZE && h_count < i_worm_x[5015:5010] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5015:5010] * PIXEL_SIZE && v_count < i_worm_y[5015:5010] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (836 < i_size && h_count >= i_worm_x[5021:5016] * PIXEL_SIZE && h_count < i_worm_x[5021:5016] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5021:5016] * PIXEL_SIZE && v_count < i_worm_y[5021:5016] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (837 < i_size && h_count >= i_worm_x[5027:5022] * PIXEL_SIZE && h_count < i_worm_x[5027:5022] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5027:5022] * PIXEL_SIZE && v_count < i_worm_y[5027:5022] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (838 < i_size && h_count >= i_worm_x[5033:5028] * PIXEL_SIZE && h_count < i_worm_x[5033:5028] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5033:5028] * PIXEL_SIZE && v_count < i_worm_y[5033:5028] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (839 < i_size && h_count >= i_worm_x[5039:5034] * PIXEL_SIZE && h_count < i_worm_x[5039:5034] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5039:5034] * PIXEL_SIZE && v_count < i_worm_y[5039:5034] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (840 < i_size && h_count >= i_worm_x[5045:5040] * PIXEL_SIZE && h_count < i_worm_x[5045:5040] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5045:5040] * PIXEL_SIZE && v_count < i_worm_y[5045:5040] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (841 < i_size && h_count >= i_worm_x[5051:5046] * PIXEL_SIZE && h_count < i_worm_x[5051:5046] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5051:5046] * PIXEL_SIZE && v_count < i_worm_y[5051:5046] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (842 < i_size && h_count >= i_worm_x[5057:5052] * PIXEL_SIZE && h_count < i_worm_x[5057:5052] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5057:5052] * PIXEL_SIZE && v_count < i_worm_y[5057:5052] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (843 < i_size && h_count >= i_worm_x[5063:5058] * PIXEL_SIZE && h_count < i_worm_x[5063:5058] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5063:5058] * PIXEL_SIZE && v_count < i_worm_y[5063:5058] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (844 < i_size && h_count >= i_worm_x[5069:5064] * PIXEL_SIZE && h_count < i_worm_x[5069:5064] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5069:5064] * PIXEL_SIZE && v_count < i_worm_y[5069:5064] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (845 < i_size && h_count >= i_worm_x[5075:5070] * PIXEL_SIZE && h_count < i_worm_x[5075:5070] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5075:5070] * PIXEL_SIZE && v_count < i_worm_y[5075:5070] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (846 < i_size && h_count >= i_worm_x[5081:5076] * PIXEL_SIZE && h_count < i_worm_x[5081:5076] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5081:5076] * PIXEL_SIZE && v_count < i_worm_y[5081:5076] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (847 < i_size && h_count >= i_worm_x[5087:5082] * PIXEL_SIZE && h_count < i_worm_x[5087:5082] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5087:5082] * PIXEL_SIZE && v_count < i_worm_y[5087:5082] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (848 < i_size && h_count >= i_worm_x[5093:5088] * PIXEL_SIZE && h_count < i_worm_x[5093:5088] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5093:5088] * PIXEL_SIZE && v_count < i_worm_y[5093:5088] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (849 < i_size && h_count >= i_worm_x[5099:5094] * PIXEL_SIZE && h_count < i_worm_x[5099:5094] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5099:5094] * PIXEL_SIZE && v_count < i_worm_y[5099:5094] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (850 < i_size && h_count >= i_worm_x[5105:5100] * PIXEL_SIZE && h_count < i_worm_x[5105:5100] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5105:5100] * PIXEL_SIZE && v_count < i_worm_y[5105:5100] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (851 < i_size && h_count >= i_worm_x[5111:5106] * PIXEL_SIZE && h_count < i_worm_x[5111:5106] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5111:5106] * PIXEL_SIZE && v_count < i_worm_y[5111:5106] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (852 < i_size && h_count >= i_worm_x[5117:5112] * PIXEL_SIZE && h_count < i_worm_x[5117:5112] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5117:5112] * PIXEL_SIZE && v_count < i_worm_y[5117:5112] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (853 < i_size && h_count >= i_worm_x[5123:5118] * PIXEL_SIZE && h_count < i_worm_x[5123:5118] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5123:5118] * PIXEL_SIZE && v_count < i_worm_y[5123:5118] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (854 < i_size && h_count >= i_worm_x[5129:5124] * PIXEL_SIZE && h_count < i_worm_x[5129:5124] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5129:5124] * PIXEL_SIZE && v_count < i_worm_y[5129:5124] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (855 < i_size && h_count >= i_worm_x[5135:5130] * PIXEL_SIZE && h_count < i_worm_x[5135:5130] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5135:5130] * PIXEL_SIZE && v_count < i_worm_y[5135:5130] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (856 < i_size && h_count >= i_worm_x[5141:5136] * PIXEL_SIZE && h_count < i_worm_x[5141:5136] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5141:5136] * PIXEL_SIZE && v_count < i_worm_y[5141:5136] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (857 < i_size && h_count >= i_worm_x[5147:5142] * PIXEL_SIZE && h_count < i_worm_x[5147:5142] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5147:5142] * PIXEL_SIZE && v_count < i_worm_y[5147:5142] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (858 < i_size && h_count >= i_worm_x[5153:5148] * PIXEL_SIZE && h_count < i_worm_x[5153:5148] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5153:5148] * PIXEL_SIZE && v_count < i_worm_y[5153:5148] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (859 < i_size && h_count >= i_worm_x[5159:5154] * PIXEL_SIZE && h_count < i_worm_x[5159:5154] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5159:5154] * PIXEL_SIZE && v_count < i_worm_y[5159:5154] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (860 < i_size && h_count >= i_worm_x[5165:5160] * PIXEL_SIZE && h_count < i_worm_x[5165:5160] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5165:5160] * PIXEL_SIZE && v_count < i_worm_y[5165:5160] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (861 < i_size && h_count >= i_worm_x[5171:5166] * PIXEL_SIZE && h_count < i_worm_x[5171:5166] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5171:5166] * PIXEL_SIZE && v_count < i_worm_y[5171:5166] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (862 < i_size && h_count >= i_worm_x[5177:5172] * PIXEL_SIZE && h_count < i_worm_x[5177:5172] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5177:5172] * PIXEL_SIZE && v_count < i_worm_y[5177:5172] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (863 < i_size && h_count >= i_worm_x[5183:5178] * PIXEL_SIZE && h_count < i_worm_x[5183:5178] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5183:5178] * PIXEL_SIZE && v_count < i_worm_y[5183:5178] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (864 < i_size && h_count >= i_worm_x[5189:5184] * PIXEL_SIZE && h_count < i_worm_x[5189:5184] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5189:5184] * PIXEL_SIZE && v_count < i_worm_y[5189:5184] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (865 < i_size && h_count >= i_worm_x[5195:5190] * PIXEL_SIZE && h_count < i_worm_x[5195:5190] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5195:5190] * PIXEL_SIZE && v_count < i_worm_y[5195:5190] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (866 < i_size && h_count >= i_worm_x[5201:5196] * PIXEL_SIZE && h_count < i_worm_x[5201:5196] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5201:5196] * PIXEL_SIZE && v_count < i_worm_y[5201:5196] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (867 < i_size && h_count >= i_worm_x[5207:5202] * PIXEL_SIZE && h_count < i_worm_x[5207:5202] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5207:5202] * PIXEL_SIZE && v_count < i_worm_y[5207:5202] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (868 < i_size && h_count >= i_worm_x[5213:5208] * PIXEL_SIZE && h_count < i_worm_x[5213:5208] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5213:5208] * PIXEL_SIZE && v_count < i_worm_y[5213:5208] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (869 < i_size && h_count >= i_worm_x[5219:5214] * PIXEL_SIZE && h_count < i_worm_x[5219:5214] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5219:5214] * PIXEL_SIZE && v_count < i_worm_y[5219:5214] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (870 < i_size && h_count >= i_worm_x[5225:5220] * PIXEL_SIZE && h_count < i_worm_x[5225:5220] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5225:5220] * PIXEL_SIZE && v_count < i_worm_y[5225:5220] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (871 < i_size && h_count >= i_worm_x[5231:5226] * PIXEL_SIZE && h_count < i_worm_x[5231:5226] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5231:5226] * PIXEL_SIZE && v_count < i_worm_y[5231:5226] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (872 < i_size && h_count >= i_worm_x[5237:5232] * PIXEL_SIZE && h_count < i_worm_x[5237:5232] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5237:5232] * PIXEL_SIZE && v_count < i_worm_y[5237:5232] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (873 < i_size && h_count >= i_worm_x[5243:5238] * PIXEL_SIZE && h_count < i_worm_x[5243:5238] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5243:5238] * PIXEL_SIZE && v_count < i_worm_y[5243:5238] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (874 < i_size && h_count >= i_worm_x[5249:5244] * PIXEL_SIZE && h_count < i_worm_x[5249:5244] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5249:5244] * PIXEL_SIZE && v_count < i_worm_y[5249:5244] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (875 < i_size && h_count >= i_worm_x[5255:5250] * PIXEL_SIZE && h_count < i_worm_x[5255:5250] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5255:5250] * PIXEL_SIZE && v_count < i_worm_y[5255:5250] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (876 < i_size && h_count >= i_worm_x[5261:5256] * PIXEL_SIZE && h_count < i_worm_x[5261:5256] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5261:5256] * PIXEL_SIZE && v_count < i_worm_y[5261:5256] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (877 < i_size && h_count >= i_worm_x[5267:5262] * PIXEL_SIZE && h_count < i_worm_x[5267:5262] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5267:5262] * PIXEL_SIZE && v_count < i_worm_y[5267:5262] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (878 < i_size && h_count >= i_worm_x[5273:5268] * PIXEL_SIZE && h_count < i_worm_x[5273:5268] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5273:5268] * PIXEL_SIZE && v_count < i_worm_y[5273:5268] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (879 < i_size && h_count >= i_worm_x[5279:5274] * PIXEL_SIZE && h_count < i_worm_x[5279:5274] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5279:5274] * PIXEL_SIZE && v_count < i_worm_y[5279:5274] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (880 < i_size && h_count >= i_worm_x[5285:5280] * PIXEL_SIZE && h_count < i_worm_x[5285:5280] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5285:5280] * PIXEL_SIZE && v_count < i_worm_y[5285:5280] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (881 < i_size && h_count >= i_worm_x[5291:5286] * PIXEL_SIZE && h_count < i_worm_x[5291:5286] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5291:5286] * PIXEL_SIZE && v_count < i_worm_y[5291:5286] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (882 < i_size && h_count >= i_worm_x[5297:5292] * PIXEL_SIZE && h_count < i_worm_x[5297:5292] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5297:5292] * PIXEL_SIZE && v_count < i_worm_y[5297:5292] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (883 < i_size && h_count >= i_worm_x[5303:5298] * PIXEL_SIZE && h_count < i_worm_x[5303:5298] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5303:5298] * PIXEL_SIZE && v_count < i_worm_y[5303:5298] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (884 < i_size && h_count >= i_worm_x[5309:5304] * PIXEL_SIZE && h_count < i_worm_x[5309:5304] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5309:5304] * PIXEL_SIZE && v_count < i_worm_y[5309:5304] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (885 < i_size && h_count >= i_worm_x[5315:5310] * PIXEL_SIZE && h_count < i_worm_x[5315:5310] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5315:5310] * PIXEL_SIZE && v_count < i_worm_y[5315:5310] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (886 < i_size && h_count >= i_worm_x[5321:5316] * PIXEL_SIZE && h_count < i_worm_x[5321:5316] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5321:5316] * PIXEL_SIZE && v_count < i_worm_y[5321:5316] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (887 < i_size && h_count >= i_worm_x[5327:5322] * PIXEL_SIZE && h_count < i_worm_x[5327:5322] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5327:5322] * PIXEL_SIZE && v_count < i_worm_y[5327:5322] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (888 < i_size && h_count >= i_worm_x[5333:5328] * PIXEL_SIZE && h_count < i_worm_x[5333:5328] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5333:5328] * PIXEL_SIZE && v_count < i_worm_y[5333:5328] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (889 < i_size && h_count >= i_worm_x[5339:5334] * PIXEL_SIZE && h_count < i_worm_x[5339:5334] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5339:5334] * PIXEL_SIZE && v_count < i_worm_y[5339:5334] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (890 < i_size && h_count >= i_worm_x[5345:5340] * PIXEL_SIZE && h_count < i_worm_x[5345:5340] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5345:5340] * PIXEL_SIZE && v_count < i_worm_y[5345:5340] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (891 < i_size && h_count >= i_worm_x[5351:5346] * PIXEL_SIZE && h_count < i_worm_x[5351:5346] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5351:5346] * PIXEL_SIZE && v_count < i_worm_y[5351:5346] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (892 < i_size && h_count >= i_worm_x[5357:5352] * PIXEL_SIZE && h_count < i_worm_x[5357:5352] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5357:5352] * PIXEL_SIZE && v_count < i_worm_y[5357:5352] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (893 < i_size && h_count >= i_worm_x[5363:5358] * PIXEL_SIZE && h_count < i_worm_x[5363:5358] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5363:5358] * PIXEL_SIZE && v_count < i_worm_y[5363:5358] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (894 < i_size && h_count >= i_worm_x[5369:5364] * PIXEL_SIZE && h_count < i_worm_x[5369:5364] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5369:5364] * PIXEL_SIZE && v_count < i_worm_y[5369:5364] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (895 < i_size && h_count >= i_worm_x[5375:5370] * PIXEL_SIZE && h_count < i_worm_x[5375:5370] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5375:5370] * PIXEL_SIZE && v_count < i_worm_y[5375:5370] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (896 < i_size && h_count >= i_worm_x[5381:5376] * PIXEL_SIZE && h_count < i_worm_x[5381:5376] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5381:5376] * PIXEL_SIZE && v_count < i_worm_y[5381:5376] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (897 < i_size && h_count >= i_worm_x[5387:5382] * PIXEL_SIZE && h_count < i_worm_x[5387:5382] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5387:5382] * PIXEL_SIZE && v_count < i_worm_y[5387:5382] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (898 < i_size && h_count >= i_worm_x[5393:5388] * PIXEL_SIZE && h_count < i_worm_x[5393:5388] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5393:5388] * PIXEL_SIZE && v_count < i_worm_y[5393:5388] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (899 < i_size && h_count >= i_worm_x[5399:5394] * PIXEL_SIZE && h_count < i_worm_x[5399:5394] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5399:5394] * PIXEL_SIZE && v_count < i_worm_y[5399:5394] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (900 < i_size && h_count >= i_worm_x[5405:5400] * PIXEL_SIZE && h_count < i_worm_x[5405:5400] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5405:5400] * PIXEL_SIZE && v_count < i_worm_y[5405:5400] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (901 < i_size && h_count >= i_worm_x[5411:5406] * PIXEL_SIZE && h_count < i_worm_x[5411:5406] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5411:5406] * PIXEL_SIZE && v_count < i_worm_y[5411:5406] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (902 < i_size && h_count >= i_worm_x[5417:5412] * PIXEL_SIZE && h_count < i_worm_x[5417:5412] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5417:5412] * PIXEL_SIZE && v_count < i_worm_y[5417:5412] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (903 < i_size && h_count >= i_worm_x[5423:5418] * PIXEL_SIZE && h_count < i_worm_x[5423:5418] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5423:5418] * PIXEL_SIZE && v_count < i_worm_y[5423:5418] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (904 < i_size && h_count >= i_worm_x[5429:5424] * PIXEL_SIZE && h_count < i_worm_x[5429:5424] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5429:5424] * PIXEL_SIZE && v_count < i_worm_y[5429:5424] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (905 < i_size && h_count >= i_worm_x[5435:5430] * PIXEL_SIZE && h_count < i_worm_x[5435:5430] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5435:5430] * PIXEL_SIZE && v_count < i_worm_y[5435:5430] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (906 < i_size && h_count >= i_worm_x[5441:5436] * PIXEL_SIZE && h_count < i_worm_x[5441:5436] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5441:5436] * PIXEL_SIZE && v_count < i_worm_y[5441:5436] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (907 < i_size && h_count >= i_worm_x[5447:5442] * PIXEL_SIZE && h_count < i_worm_x[5447:5442] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5447:5442] * PIXEL_SIZE && v_count < i_worm_y[5447:5442] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (908 < i_size && h_count >= i_worm_x[5453:5448] * PIXEL_SIZE && h_count < i_worm_x[5453:5448] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5453:5448] * PIXEL_SIZE && v_count < i_worm_y[5453:5448] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (909 < i_size && h_count >= i_worm_x[5459:5454] * PIXEL_SIZE && h_count < i_worm_x[5459:5454] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5459:5454] * PIXEL_SIZE && v_count < i_worm_y[5459:5454] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (910 < i_size && h_count >= i_worm_x[5465:5460] * PIXEL_SIZE && h_count < i_worm_x[5465:5460] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5465:5460] * PIXEL_SIZE && v_count < i_worm_y[5465:5460] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (911 < i_size && h_count >= i_worm_x[5471:5466] * PIXEL_SIZE && h_count < i_worm_x[5471:5466] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5471:5466] * PIXEL_SIZE && v_count < i_worm_y[5471:5466] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (912 < i_size && h_count >= i_worm_x[5477:5472] * PIXEL_SIZE && h_count < i_worm_x[5477:5472] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5477:5472] * PIXEL_SIZE && v_count < i_worm_y[5477:5472] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (913 < i_size && h_count >= i_worm_x[5483:5478] * PIXEL_SIZE && h_count < i_worm_x[5483:5478] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5483:5478] * PIXEL_SIZE && v_count < i_worm_y[5483:5478] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (914 < i_size && h_count >= i_worm_x[5489:5484] * PIXEL_SIZE && h_count < i_worm_x[5489:5484] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5489:5484] * PIXEL_SIZE && v_count < i_worm_y[5489:5484] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (915 < i_size && h_count >= i_worm_x[5495:5490] * PIXEL_SIZE && h_count < i_worm_x[5495:5490] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5495:5490] * PIXEL_SIZE && v_count < i_worm_y[5495:5490] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (916 < i_size && h_count >= i_worm_x[5501:5496] * PIXEL_SIZE && h_count < i_worm_x[5501:5496] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5501:5496] * PIXEL_SIZE && v_count < i_worm_y[5501:5496] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (917 < i_size && h_count >= i_worm_x[5507:5502] * PIXEL_SIZE && h_count < i_worm_x[5507:5502] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5507:5502] * PIXEL_SIZE && v_count < i_worm_y[5507:5502] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (918 < i_size && h_count >= i_worm_x[5513:5508] * PIXEL_SIZE && h_count < i_worm_x[5513:5508] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5513:5508] * PIXEL_SIZE && v_count < i_worm_y[5513:5508] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (919 < i_size && h_count >= i_worm_x[5519:5514] * PIXEL_SIZE && h_count < i_worm_x[5519:5514] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5519:5514] * PIXEL_SIZE && v_count < i_worm_y[5519:5514] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (920 < i_size && h_count >= i_worm_x[5525:5520] * PIXEL_SIZE && h_count < i_worm_x[5525:5520] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5525:5520] * PIXEL_SIZE && v_count < i_worm_y[5525:5520] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (921 < i_size && h_count >= i_worm_x[5531:5526] * PIXEL_SIZE && h_count < i_worm_x[5531:5526] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5531:5526] * PIXEL_SIZE && v_count < i_worm_y[5531:5526] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (922 < i_size && h_count >= i_worm_x[5537:5532] * PIXEL_SIZE && h_count < i_worm_x[5537:5532] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5537:5532] * PIXEL_SIZE && v_count < i_worm_y[5537:5532] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (923 < i_size && h_count >= i_worm_x[5543:5538] * PIXEL_SIZE && h_count < i_worm_x[5543:5538] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5543:5538] * PIXEL_SIZE && v_count < i_worm_y[5543:5538] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (924 < i_size && h_count >= i_worm_x[5549:5544] * PIXEL_SIZE && h_count < i_worm_x[5549:5544] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5549:5544] * PIXEL_SIZE && v_count < i_worm_y[5549:5544] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (925 < i_size && h_count >= i_worm_x[5555:5550] * PIXEL_SIZE && h_count < i_worm_x[5555:5550] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5555:5550] * PIXEL_SIZE && v_count < i_worm_y[5555:5550] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (926 < i_size && h_count >= i_worm_x[5561:5556] * PIXEL_SIZE && h_count < i_worm_x[5561:5556] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5561:5556] * PIXEL_SIZE && v_count < i_worm_y[5561:5556] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (927 < i_size && h_count >= i_worm_x[5567:5562] * PIXEL_SIZE && h_count < i_worm_x[5567:5562] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5567:5562] * PIXEL_SIZE && v_count < i_worm_y[5567:5562] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (928 < i_size && h_count >= i_worm_x[5573:5568] * PIXEL_SIZE && h_count < i_worm_x[5573:5568] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5573:5568] * PIXEL_SIZE && v_count < i_worm_y[5573:5568] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (929 < i_size && h_count >= i_worm_x[5579:5574] * PIXEL_SIZE && h_count < i_worm_x[5579:5574] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5579:5574] * PIXEL_SIZE && v_count < i_worm_y[5579:5574] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (930 < i_size && h_count >= i_worm_x[5585:5580] * PIXEL_SIZE && h_count < i_worm_x[5585:5580] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5585:5580] * PIXEL_SIZE && v_count < i_worm_y[5585:5580] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (931 < i_size && h_count >= i_worm_x[5591:5586] * PIXEL_SIZE && h_count < i_worm_x[5591:5586] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5591:5586] * PIXEL_SIZE && v_count < i_worm_y[5591:5586] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (932 < i_size && h_count >= i_worm_x[5597:5592] * PIXEL_SIZE && h_count < i_worm_x[5597:5592] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5597:5592] * PIXEL_SIZE && v_count < i_worm_y[5597:5592] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (933 < i_size && h_count >= i_worm_x[5603:5598] * PIXEL_SIZE && h_count < i_worm_x[5603:5598] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5603:5598] * PIXEL_SIZE && v_count < i_worm_y[5603:5598] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (934 < i_size && h_count >= i_worm_x[5609:5604] * PIXEL_SIZE && h_count < i_worm_x[5609:5604] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5609:5604] * PIXEL_SIZE && v_count < i_worm_y[5609:5604] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (935 < i_size && h_count >= i_worm_x[5615:5610] * PIXEL_SIZE && h_count < i_worm_x[5615:5610] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5615:5610] * PIXEL_SIZE && v_count < i_worm_y[5615:5610] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (936 < i_size && h_count >= i_worm_x[5621:5616] * PIXEL_SIZE && h_count < i_worm_x[5621:5616] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5621:5616] * PIXEL_SIZE && v_count < i_worm_y[5621:5616] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (937 < i_size && h_count >= i_worm_x[5627:5622] * PIXEL_SIZE && h_count < i_worm_x[5627:5622] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5627:5622] * PIXEL_SIZE && v_count < i_worm_y[5627:5622] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (938 < i_size && h_count >= i_worm_x[5633:5628] * PIXEL_SIZE && h_count < i_worm_x[5633:5628] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5633:5628] * PIXEL_SIZE && v_count < i_worm_y[5633:5628] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (939 < i_size && h_count >= i_worm_x[5639:5634] * PIXEL_SIZE && h_count < i_worm_x[5639:5634] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5639:5634] * PIXEL_SIZE && v_count < i_worm_y[5639:5634] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (940 < i_size && h_count >= i_worm_x[5645:5640] * PIXEL_SIZE && h_count < i_worm_x[5645:5640] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5645:5640] * PIXEL_SIZE && v_count < i_worm_y[5645:5640] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (941 < i_size && h_count >= i_worm_x[5651:5646] * PIXEL_SIZE && h_count < i_worm_x[5651:5646] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5651:5646] * PIXEL_SIZE && v_count < i_worm_y[5651:5646] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (942 < i_size && h_count >= i_worm_x[5657:5652] * PIXEL_SIZE && h_count < i_worm_x[5657:5652] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5657:5652] * PIXEL_SIZE && v_count < i_worm_y[5657:5652] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (943 < i_size && h_count >= i_worm_x[5663:5658] * PIXEL_SIZE && h_count < i_worm_x[5663:5658] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5663:5658] * PIXEL_SIZE && v_count < i_worm_y[5663:5658] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (944 < i_size && h_count >= i_worm_x[5669:5664] * PIXEL_SIZE && h_count < i_worm_x[5669:5664] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5669:5664] * PIXEL_SIZE && v_count < i_worm_y[5669:5664] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (945 < i_size && h_count >= i_worm_x[5675:5670] * PIXEL_SIZE && h_count < i_worm_x[5675:5670] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5675:5670] * PIXEL_SIZE && v_count < i_worm_y[5675:5670] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (946 < i_size && h_count >= i_worm_x[5681:5676] * PIXEL_SIZE && h_count < i_worm_x[5681:5676] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5681:5676] * PIXEL_SIZE && v_count < i_worm_y[5681:5676] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (947 < i_size && h_count >= i_worm_x[5687:5682] * PIXEL_SIZE && h_count < i_worm_x[5687:5682] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5687:5682] * PIXEL_SIZE && v_count < i_worm_y[5687:5682] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (948 < i_size && h_count >= i_worm_x[5693:5688] * PIXEL_SIZE && h_count < i_worm_x[5693:5688] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5693:5688] * PIXEL_SIZE && v_count < i_worm_y[5693:5688] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (949 < i_size && h_count >= i_worm_x[5699:5694] * PIXEL_SIZE && h_count < i_worm_x[5699:5694] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5699:5694] * PIXEL_SIZE && v_count < i_worm_y[5699:5694] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (950 < i_size && h_count >= i_worm_x[5705:5700] * PIXEL_SIZE && h_count < i_worm_x[5705:5700] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5705:5700] * PIXEL_SIZE && v_count < i_worm_y[5705:5700] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (951 < i_size && h_count >= i_worm_x[5711:5706] * PIXEL_SIZE && h_count < i_worm_x[5711:5706] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5711:5706] * PIXEL_SIZE && v_count < i_worm_y[5711:5706] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (952 < i_size && h_count >= i_worm_x[5717:5712] * PIXEL_SIZE && h_count < i_worm_x[5717:5712] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5717:5712] * PIXEL_SIZE && v_count < i_worm_y[5717:5712] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (953 < i_size && h_count >= i_worm_x[5723:5718] * PIXEL_SIZE && h_count < i_worm_x[5723:5718] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5723:5718] * PIXEL_SIZE && v_count < i_worm_y[5723:5718] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (954 < i_size && h_count >= i_worm_x[5729:5724] * PIXEL_SIZE && h_count < i_worm_x[5729:5724] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5729:5724] * PIXEL_SIZE && v_count < i_worm_y[5729:5724] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (955 < i_size && h_count >= i_worm_x[5735:5730] * PIXEL_SIZE && h_count < i_worm_x[5735:5730] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5735:5730] * PIXEL_SIZE && v_count < i_worm_y[5735:5730] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (956 < i_size && h_count >= i_worm_x[5741:5736] * PIXEL_SIZE && h_count < i_worm_x[5741:5736] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5741:5736] * PIXEL_SIZE && v_count < i_worm_y[5741:5736] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (957 < i_size && h_count >= i_worm_x[5747:5742] * PIXEL_SIZE && h_count < i_worm_x[5747:5742] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5747:5742] * PIXEL_SIZE && v_count < i_worm_y[5747:5742] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (958 < i_size && h_count >= i_worm_x[5753:5748] * PIXEL_SIZE && h_count < i_worm_x[5753:5748] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5753:5748] * PIXEL_SIZE && v_count < i_worm_y[5753:5748] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (959 < i_size && h_count >= i_worm_x[5759:5754] * PIXEL_SIZE && h_count < i_worm_x[5759:5754] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5759:5754] * PIXEL_SIZE && v_count < i_worm_y[5759:5754] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (960 < i_size && h_count >= i_worm_x[5765:5760] * PIXEL_SIZE && h_count < i_worm_x[5765:5760] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5765:5760] * PIXEL_SIZE && v_count < i_worm_y[5765:5760] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (961 < i_size && h_count >= i_worm_x[5771:5766] * PIXEL_SIZE && h_count < i_worm_x[5771:5766] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5771:5766] * PIXEL_SIZE && v_count < i_worm_y[5771:5766] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (962 < i_size && h_count >= i_worm_x[5777:5772] * PIXEL_SIZE && h_count < i_worm_x[5777:5772] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5777:5772] * PIXEL_SIZE && v_count < i_worm_y[5777:5772] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (963 < i_size && h_count >= i_worm_x[5783:5778] * PIXEL_SIZE && h_count < i_worm_x[5783:5778] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5783:5778] * PIXEL_SIZE && v_count < i_worm_y[5783:5778] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (964 < i_size && h_count >= i_worm_x[5789:5784] * PIXEL_SIZE && h_count < i_worm_x[5789:5784] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5789:5784] * PIXEL_SIZE && v_count < i_worm_y[5789:5784] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (965 < i_size && h_count >= i_worm_x[5795:5790] * PIXEL_SIZE && h_count < i_worm_x[5795:5790] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5795:5790] * PIXEL_SIZE && v_count < i_worm_y[5795:5790] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (966 < i_size && h_count >= i_worm_x[5801:5796] * PIXEL_SIZE && h_count < i_worm_x[5801:5796] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5801:5796] * PIXEL_SIZE && v_count < i_worm_y[5801:5796] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (967 < i_size && h_count >= i_worm_x[5807:5802] * PIXEL_SIZE && h_count < i_worm_x[5807:5802] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5807:5802] * PIXEL_SIZE && v_count < i_worm_y[5807:5802] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (968 < i_size && h_count >= i_worm_x[5813:5808] * PIXEL_SIZE && h_count < i_worm_x[5813:5808] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5813:5808] * PIXEL_SIZE && v_count < i_worm_y[5813:5808] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (969 < i_size && h_count >= i_worm_x[5819:5814] * PIXEL_SIZE && h_count < i_worm_x[5819:5814] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5819:5814] * PIXEL_SIZE && v_count < i_worm_y[5819:5814] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (970 < i_size && h_count >= i_worm_x[5825:5820] * PIXEL_SIZE && h_count < i_worm_x[5825:5820] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5825:5820] * PIXEL_SIZE && v_count < i_worm_y[5825:5820] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (971 < i_size && h_count >= i_worm_x[5831:5826] * PIXEL_SIZE && h_count < i_worm_x[5831:5826] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5831:5826] * PIXEL_SIZE && v_count < i_worm_y[5831:5826] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (972 < i_size && h_count >= i_worm_x[5837:5832] * PIXEL_SIZE && h_count < i_worm_x[5837:5832] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5837:5832] * PIXEL_SIZE && v_count < i_worm_y[5837:5832] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (973 < i_size && h_count >= i_worm_x[5843:5838] * PIXEL_SIZE && h_count < i_worm_x[5843:5838] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5843:5838] * PIXEL_SIZE && v_count < i_worm_y[5843:5838] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (974 < i_size && h_count >= i_worm_x[5849:5844] * PIXEL_SIZE && h_count < i_worm_x[5849:5844] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5849:5844] * PIXEL_SIZE && v_count < i_worm_y[5849:5844] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (975 < i_size && h_count >= i_worm_x[5855:5850] * PIXEL_SIZE && h_count < i_worm_x[5855:5850] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5855:5850] * PIXEL_SIZE && v_count < i_worm_y[5855:5850] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (976 < i_size && h_count >= i_worm_x[5861:5856] * PIXEL_SIZE && h_count < i_worm_x[5861:5856] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5861:5856] * PIXEL_SIZE && v_count < i_worm_y[5861:5856] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (977 < i_size && h_count >= i_worm_x[5867:5862] * PIXEL_SIZE && h_count < i_worm_x[5867:5862] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5867:5862] * PIXEL_SIZE && v_count < i_worm_y[5867:5862] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (978 < i_size && h_count >= i_worm_x[5873:5868] * PIXEL_SIZE && h_count < i_worm_x[5873:5868] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5873:5868] * PIXEL_SIZE && v_count < i_worm_y[5873:5868] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (979 < i_size && h_count >= i_worm_x[5879:5874] * PIXEL_SIZE && h_count < i_worm_x[5879:5874] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5879:5874] * PIXEL_SIZE && v_count < i_worm_y[5879:5874] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (980 < i_size && h_count >= i_worm_x[5885:5880] * PIXEL_SIZE && h_count < i_worm_x[5885:5880] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5885:5880] * PIXEL_SIZE && v_count < i_worm_y[5885:5880] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (981 < i_size && h_count >= i_worm_x[5891:5886] * PIXEL_SIZE && h_count < i_worm_x[5891:5886] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5891:5886] * PIXEL_SIZE && v_count < i_worm_y[5891:5886] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (982 < i_size && h_count >= i_worm_x[5897:5892] * PIXEL_SIZE && h_count < i_worm_x[5897:5892] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5897:5892] * PIXEL_SIZE && v_count < i_worm_y[5897:5892] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (983 < i_size && h_count >= i_worm_x[5903:5898] * PIXEL_SIZE && h_count < i_worm_x[5903:5898] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5903:5898] * PIXEL_SIZE && v_count < i_worm_y[5903:5898] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (984 < i_size && h_count >= i_worm_x[5909:5904] * PIXEL_SIZE && h_count < i_worm_x[5909:5904] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5909:5904] * PIXEL_SIZE && v_count < i_worm_y[5909:5904] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (985 < i_size && h_count >= i_worm_x[5915:5910] * PIXEL_SIZE && h_count < i_worm_x[5915:5910] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5915:5910] * PIXEL_SIZE && v_count < i_worm_y[5915:5910] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (986 < i_size && h_count >= i_worm_x[5921:5916] * PIXEL_SIZE && h_count < i_worm_x[5921:5916] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5921:5916] * PIXEL_SIZE && v_count < i_worm_y[5921:5916] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (987 < i_size && h_count >= i_worm_x[5927:5922] * PIXEL_SIZE && h_count < i_worm_x[5927:5922] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5927:5922] * PIXEL_SIZE && v_count < i_worm_y[5927:5922] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (988 < i_size && h_count >= i_worm_x[5933:5928] * PIXEL_SIZE && h_count < i_worm_x[5933:5928] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5933:5928] * PIXEL_SIZE && v_count < i_worm_y[5933:5928] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (989 < i_size && h_count >= i_worm_x[5939:5934] * PIXEL_SIZE && h_count < i_worm_x[5939:5934] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5939:5934] * PIXEL_SIZE && v_count < i_worm_y[5939:5934] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (990 < i_size && h_count >= i_worm_x[5945:5940] * PIXEL_SIZE && h_count < i_worm_x[5945:5940] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5945:5940] * PIXEL_SIZE && v_count < i_worm_y[5945:5940] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (991 < i_size && h_count >= i_worm_x[5951:5946] * PIXEL_SIZE && h_count < i_worm_x[5951:5946] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5951:5946] * PIXEL_SIZE && v_count < i_worm_y[5951:5946] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (992 < i_size && h_count >= i_worm_x[5957:5952] * PIXEL_SIZE && h_count < i_worm_x[5957:5952] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5957:5952] * PIXEL_SIZE && v_count < i_worm_y[5957:5952] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (993 < i_size && h_count >= i_worm_x[5963:5958] * PIXEL_SIZE && h_count < i_worm_x[5963:5958] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5963:5958] * PIXEL_SIZE && v_count < i_worm_y[5963:5958] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (994 < i_size && h_count >= i_worm_x[5969:5964] * PIXEL_SIZE && h_count < i_worm_x[5969:5964] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5969:5964] * PIXEL_SIZE && v_count < i_worm_y[5969:5964] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (995 < i_size && h_count >= i_worm_x[5975:5970] * PIXEL_SIZE && h_count < i_worm_x[5975:5970] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5975:5970] * PIXEL_SIZE && v_count < i_worm_y[5975:5970] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (996 < i_size && h_count >= i_worm_x[5981:5976] * PIXEL_SIZE && h_count < i_worm_x[5981:5976] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5981:5976] * PIXEL_SIZE && v_count < i_worm_y[5981:5976] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (997 < i_size && h_count >= i_worm_x[5987:5982] * PIXEL_SIZE && h_count < i_worm_x[5987:5982] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5987:5982] * PIXEL_SIZE && v_count < i_worm_y[5987:5982] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (998 < i_size && h_count >= i_worm_x[5993:5988] * PIXEL_SIZE && h_count < i_worm_x[5993:5988] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5993:5988] * PIXEL_SIZE && v_count < i_worm_y[5993:5988] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (999 < i_size && h_count >= i_worm_x[5999:5994] * PIXEL_SIZE && h_count < i_worm_x[5999:5994] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[5999:5994] * PIXEL_SIZE && v_count < i_worm_y[5999:5994] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1000 < i_size && h_count >= i_worm_x[6005:6000] * PIXEL_SIZE && h_count < i_worm_x[6005:6000] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6005:6000] * PIXEL_SIZE && v_count < i_worm_y[6005:6000] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1001 < i_size && h_count >= i_worm_x[6011:6006] * PIXEL_SIZE && h_count < i_worm_x[6011:6006] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6011:6006] * PIXEL_SIZE && v_count < i_worm_y[6011:6006] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1002 < i_size && h_count >= i_worm_x[6017:6012] * PIXEL_SIZE && h_count < i_worm_x[6017:6012] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6017:6012] * PIXEL_SIZE && v_count < i_worm_y[6017:6012] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1003 < i_size && h_count >= i_worm_x[6023:6018] * PIXEL_SIZE && h_count < i_worm_x[6023:6018] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6023:6018] * PIXEL_SIZE && v_count < i_worm_y[6023:6018] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1004 < i_size && h_count >= i_worm_x[6029:6024] * PIXEL_SIZE && h_count < i_worm_x[6029:6024] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6029:6024] * PIXEL_SIZE && v_count < i_worm_y[6029:6024] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1005 < i_size && h_count >= i_worm_x[6035:6030] * PIXEL_SIZE && h_count < i_worm_x[6035:6030] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6035:6030] * PIXEL_SIZE && v_count < i_worm_y[6035:6030] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1006 < i_size && h_count >= i_worm_x[6041:6036] * PIXEL_SIZE && h_count < i_worm_x[6041:6036] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6041:6036] * PIXEL_SIZE && v_count < i_worm_y[6041:6036] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1007 < i_size && h_count >= i_worm_x[6047:6042] * PIXEL_SIZE && h_count < i_worm_x[6047:6042] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6047:6042] * PIXEL_SIZE && v_count < i_worm_y[6047:6042] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1008 < i_size && h_count >= i_worm_x[6053:6048] * PIXEL_SIZE && h_count < i_worm_x[6053:6048] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6053:6048] * PIXEL_SIZE && v_count < i_worm_y[6053:6048] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1009 < i_size && h_count >= i_worm_x[6059:6054] * PIXEL_SIZE && h_count < i_worm_x[6059:6054] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6059:6054] * PIXEL_SIZE && v_count < i_worm_y[6059:6054] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1010 < i_size && h_count >= i_worm_x[6065:6060] * PIXEL_SIZE && h_count < i_worm_x[6065:6060] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6065:6060] * PIXEL_SIZE && v_count < i_worm_y[6065:6060] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1011 < i_size && h_count >= i_worm_x[6071:6066] * PIXEL_SIZE && h_count < i_worm_x[6071:6066] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6071:6066] * PIXEL_SIZE && v_count < i_worm_y[6071:6066] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1012 < i_size && h_count >= i_worm_x[6077:6072] * PIXEL_SIZE && h_count < i_worm_x[6077:6072] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6077:6072] * PIXEL_SIZE && v_count < i_worm_y[6077:6072] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1013 < i_size && h_count >= i_worm_x[6083:6078] * PIXEL_SIZE && h_count < i_worm_x[6083:6078] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6083:6078] * PIXEL_SIZE && v_count < i_worm_y[6083:6078] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1014 < i_size && h_count >= i_worm_x[6089:6084] * PIXEL_SIZE && h_count < i_worm_x[6089:6084] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6089:6084] * PIXEL_SIZE && v_count < i_worm_y[6089:6084] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1015 < i_size && h_count >= i_worm_x[6095:6090] * PIXEL_SIZE && h_count < i_worm_x[6095:6090] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6095:6090] * PIXEL_SIZE && v_count < i_worm_y[6095:6090] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1016 < i_size && h_count >= i_worm_x[6101:6096] * PIXEL_SIZE && h_count < i_worm_x[6101:6096] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6101:6096] * PIXEL_SIZE && v_count < i_worm_y[6101:6096] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1017 < i_size && h_count >= i_worm_x[6107:6102] * PIXEL_SIZE && h_count < i_worm_x[6107:6102] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6107:6102] * PIXEL_SIZE && v_count < i_worm_y[6107:6102] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1018 < i_size && h_count >= i_worm_x[6113:6108] * PIXEL_SIZE && h_count < i_worm_x[6113:6108] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6113:6108] * PIXEL_SIZE && v_count < i_worm_y[6113:6108] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1019 < i_size && h_count >= i_worm_x[6119:6114] * PIXEL_SIZE && h_count < i_worm_x[6119:6114] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6119:6114] * PIXEL_SIZE && v_count < i_worm_y[6119:6114] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1020 < i_size && h_count >= i_worm_x[6125:6120] * PIXEL_SIZE && h_count < i_worm_x[6125:6120] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6125:6120] * PIXEL_SIZE && v_count < i_worm_y[6125:6120] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1021 < i_size && h_count >= i_worm_x[6131:6126] * PIXEL_SIZE && h_count < i_worm_x[6131:6126] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6131:6126] * PIXEL_SIZE && v_count < i_worm_y[6131:6126] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1022 < i_size && h_count >= i_worm_x[6137:6132] * PIXEL_SIZE && h_count < i_worm_x[6137:6132] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6137:6132] * PIXEL_SIZE && v_count < i_worm_y[6137:6132] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1023 < i_size && h_count >= i_worm_x[6143:6138] * PIXEL_SIZE && h_count < i_worm_x[6143:6138] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6143:6138] * PIXEL_SIZE && v_count < i_worm_y[6143:6138] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1024 < i_size && h_count >= i_worm_x[6149:6144] * PIXEL_SIZE && h_count < i_worm_x[6149:6144] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6149:6144] * PIXEL_SIZE && v_count < i_worm_y[6149:6144] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1025 < i_size && h_count >= i_worm_x[6155:6150] * PIXEL_SIZE && h_count < i_worm_x[6155:6150] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6155:6150] * PIXEL_SIZE && v_count < i_worm_y[6155:6150] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1026 < i_size && h_count >= i_worm_x[6161:6156] * PIXEL_SIZE && h_count < i_worm_x[6161:6156] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6161:6156] * PIXEL_SIZE && v_count < i_worm_y[6161:6156] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1027 < i_size && h_count >= i_worm_x[6167:6162] * PIXEL_SIZE && h_count < i_worm_x[6167:6162] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6167:6162] * PIXEL_SIZE && v_count < i_worm_y[6167:6162] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1028 < i_size && h_count >= i_worm_x[6173:6168] * PIXEL_SIZE && h_count < i_worm_x[6173:6168] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6173:6168] * PIXEL_SIZE && v_count < i_worm_y[6173:6168] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1029 < i_size && h_count >= i_worm_x[6179:6174] * PIXEL_SIZE && h_count < i_worm_x[6179:6174] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6179:6174] * PIXEL_SIZE && v_count < i_worm_y[6179:6174] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1030 < i_size && h_count >= i_worm_x[6185:6180] * PIXEL_SIZE && h_count < i_worm_x[6185:6180] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6185:6180] * PIXEL_SIZE && v_count < i_worm_y[6185:6180] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1031 < i_size && h_count >= i_worm_x[6191:6186] * PIXEL_SIZE && h_count < i_worm_x[6191:6186] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6191:6186] * PIXEL_SIZE && v_count < i_worm_y[6191:6186] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1032 < i_size && h_count >= i_worm_x[6197:6192] * PIXEL_SIZE && h_count < i_worm_x[6197:6192] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6197:6192] * PIXEL_SIZE && v_count < i_worm_y[6197:6192] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1033 < i_size && h_count >= i_worm_x[6203:6198] * PIXEL_SIZE && h_count < i_worm_x[6203:6198] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6203:6198] * PIXEL_SIZE && v_count < i_worm_y[6203:6198] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1034 < i_size && h_count >= i_worm_x[6209:6204] * PIXEL_SIZE && h_count < i_worm_x[6209:6204] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6209:6204] * PIXEL_SIZE && v_count < i_worm_y[6209:6204] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1035 < i_size && h_count >= i_worm_x[6215:6210] * PIXEL_SIZE && h_count < i_worm_x[6215:6210] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6215:6210] * PIXEL_SIZE && v_count < i_worm_y[6215:6210] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1036 < i_size && h_count >= i_worm_x[6221:6216] * PIXEL_SIZE && h_count < i_worm_x[6221:6216] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6221:6216] * PIXEL_SIZE && v_count < i_worm_y[6221:6216] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1037 < i_size && h_count >= i_worm_x[6227:6222] * PIXEL_SIZE && h_count < i_worm_x[6227:6222] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6227:6222] * PIXEL_SIZE && v_count < i_worm_y[6227:6222] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1038 < i_size && h_count >= i_worm_x[6233:6228] * PIXEL_SIZE && h_count < i_worm_x[6233:6228] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6233:6228] * PIXEL_SIZE && v_count < i_worm_y[6233:6228] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1039 < i_size && h_count >= i_worm_x[6239:6234] * PIXEL_SIZE && h_count < i_worm_x[6239:6234] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6239:6234] * PIXEL_SIZE && v_count < i_worm_y[6239:6234] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1040 < i_size && h_count >= i_worm_x[6245:6240] * PIXEL_SIZE && h_count < i_worm_x[6245:6240] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6245:6240] * PIXEL_SIZE && v_count < i_worm_y[6245:6240] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1041 < i_size && h_count >= i_worm_x[6251:6246] * PIXEL_SIZE && h_count < i_worm_x[6251:6246] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6251:6246] * PIXEL_SIZE && v_count < i_worm_y[6251:6246] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1042 < i_size && h_count >= i_worm_x[6257:6252] * PIXEL_SIZE && h_count < i_worm_x[6257:6252] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6257:6252] * PIXEL_SIZE && v_count < i_worm_y[6257:6252] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1043 < i_size && h_count >= i_worm_x[6263:6258] * PIXEL_SIZE && h_count < i_worm_x[6263:6258] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6263:6258] * PIXEL_SIZE && v_count < i_worm_y[6263:6258] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1044 < i_size && h_count >= i_worm_x[6269:6264] * PIXEL_SIZE && h_count < i_worm_x[6269:6264] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6269:6264] * PIXEL_SIZE && v_count < i_worm_y[6269:6264] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1045 < i_size && h_count >= i_worm_x[6275:6270] * PIXEL_SIZE && h_count < i_worm_x[6275:6270] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6275:6270] * PIXEL_SIZE && v_count < i_worm_y[6275:6270] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1046 < i_size && h_count >= i_worm_x[6281:6276] * PIXEL_SIZE && h_count < i_worm_x[6281:6276] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6281:6276] * PIXEL_SIZE && v_count < i_worm_y[6281:6276] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1047 < i_size && h_count >= i_worm_x[6287:6282] * PIXEL_SIZE && h_count < i_worm_x[6287:6282] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6287:6282] * PIXEL_SIZE && v_count < i_worm_y[6287:6282] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1048 < i_size && h_count >= i_worm_x[6293:6288] * PIXEL_SIZE && h_count < i_worm_x[6293:6288] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6293:6288] * PIXEL_SIZE && v_count < i_worm_y[6293:6288] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1049 < i_size && h_count >= i_worm_x[6299:6294] * PIXEL_SIZE && h_count < i_worm_x[6299:6294] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6299:6294] * PIXEL_SIZE && v_count < i_worm_y[6299:6294] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1050 < i_size && h_count >= i_worm_x[6305:6300] * PIXEL_SIZE && h_count < i_worm_x[6305:6300] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6305:6300] * PIXEL_SIZE && v_count < i_worm_y[6305:6300] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1051 < i_size && h_count >= i_worm_x[6311:6306] * PIXEL_SIZE && h_count < i_worm_x[6311:6306] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6311:6306] * PIXEL_SIZE && v_count < i_worm_y[6311:6306] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1052 < i_size && h_count >= i_worm_x[6317:6312] * PIXEL_SIZE && h_count < i_worm_x[6317:6312] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6317:6312] * PIXEL_SIZE && v_count < i_worm_y[6317:6312] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1053 < i_size && h_count >= i_worm_x[6323:6318] * PIXEL_SIZE && h_count < i_worm_x[6323:6318] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6323:6318] * PIXEL_SIZE && v_count < i_worm_y[6323:6318] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1054 < i_size && h_count >= i_worm_x[6329:6324] * PIXEL_SIZE && h_count < i_worm_x[6329:6324] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6329:6324] * PIXEL_SIZE && v_count < i_worm_y[6329:6324] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1055 < i_size && h_count >= i_worm_x[6335:6330] * PIXEL_SIZE && h_count < i_worm_x[6335:6330] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6335:6330] * PIXEL_SIZE && v_count < i_worm_y[6335:6330] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1056 < i_size && h_count >= i_worm_x[6341:6336] * PIXEL_SIZE && h_count < i_worm_x[6341:6336] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6341:6336] * PIXEL_SIZE && v_count < i_worm_y[6341:6336] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1057 < i_size && h_count >= i_worm_x[6347:6342] * PIXEL_SIZE && h_count < i_worm_x[6347:6342] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6347:6342] * PIXEL_SIZE && v_count < i_worm_y[6347:6342] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1058 < i_size && h_count >= i_worm_x[6353:6348] * PIXEL_SIZE && h_count < i_worm_x[6353:6348] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6353:6348] * PIXEL_SIZE && v_count < i_worm_y[6353:6348] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1059 < i_size && h_count >= i_worm_x[6359:6354] * PIXEL_SIZE && h_count < i_worm_x[6359:6354] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6359:6354] * PIXEL_SIZE && v_count < i_worm_y[6359:6354] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1060 < i_size && h_count >= i_worm_x[6365:6360] * PIXEL_SIZE && h_count < i_worm_x[6365:6360] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6365:6360] * PIXEL_SIZE && v_count < i_worm_y[6365:6360] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1061 < i_size && h_count >= i_worm_x[6371:6366] * PIXEL_SIZE && h_count < i_worm_x[6371:6366] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6371:6366] * PIXEL_SIZE && v_count < i_worm_y[6371:6366] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1062 < i_size && h_count >= i_worm_x[6377:6372] * PIXEL_SIZE && h_count < i_worm_x[6377:6372] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6377:6372] * PIXEL_SIZE && v_count < i_worm_y[6377:6372] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1063 < i_size && h_count >= i_worm_x[6383:6378] * PIXEL_SIZE && h_count < i_worm_x[6383:6378] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6383:6378] * PIXEL_SIZE && v_count < i_worm_y[6383:6378] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1064 < i_size && h_count >= i_worm_x[6389:6384] * PIXEL_SIZE && h_count < i_worm_x[6389:6384] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6389:6384] * PIXEL_SIZE && v_count < i_worm_y[6389:6384] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1065 < i_size && h_count >= i_worm_x[6395:6390] * PIXEL_SIZE && h_count < i_worm_x[6395:6390] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6395:6390] * PIXEL_SIZE && v_count < i_worm_y[6395:6390] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1066 < i_size && h_count >= i_worm_x[6401:6396] * PIXEL_SIZE && h_count < i_worm_x[6401:6396] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6401:6396] * PIXEL_SIZE && v_count < i_worm_y[6401:6396] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1067 < i_size && h_count >= i_worm_x[6407:6402] * PIXEL_SIZE && h_count < i_worm_x[6407:6402] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6407:6402] * PIXEL_SIZE && v_count < i_worm_y[6407:6402] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1068 < i_size && h_count >= i_worm_x[6413:6408] * PIXEL_SIZE && h_count < i_worm_x[6413:6408] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6413:6408] * PIXEL_SIZE && v_count < i_worm_y[6413:6408] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1069 < i_size && h_count >= i_worm_x[6419:6414] * PIXEL_SIZE && h_count < i_worm_x[6419:6414] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6419:6414] * PIXEL_SIZE && v_count < i_worm_y[6419:6414] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1070 < i_size && h_count >= i_worm_x[6425:6420] * PIXEL_SIZE && h_count < i_worm_x[6425:6420] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6425:6420] * PIXEL_SIZE && v_count < i_worm_y[6425:6420] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1071 < i_size && h_count >= i_worm_x[6431:6426] * PIXEL_SIZE && h_count < i_worm_x[6431:6426] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6431:6426] * PIXEL_SIZE && v_count < i_worm_y[6431:6426] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1072 < i_size && h_count >= i_worm_x[6437:6432] * PIXEL_SIZE && h_count < i_worm_x[6437:6432] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6437:6432] * PIXEL_SIZE && v_count < i_worm_y[6437:6432] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1073 < i_size && h_count >= i_worm_x[6443:6438] * PIXEL_SIZE && h_count < i_worm_x[6443:6438] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6443:6438] * PIXEL_SIZE && v_count < i_worm_y[6443:6438] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1074 < i_size && h_count >= i_worm_x[6449:6444] * PIXEL_SIZE && h_count < i_worm_x[6449:6444] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6449:6444] * PIXEL_SIZE && v_count < i_worm_y[6449:6444] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1075 < i_size && h_count >= i_worm_x[6455:6450] * PIXEL_SIZE && h_count < i_worm_x[6455:6450] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6455:6450] * PIXEL_SIZE && v_count < i_worm_y[6455:6450] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1076 < i_size && h_count >= i_worm_x[6461:6456] * PIXEL_SIZE && h_count < i_worm_x[6461:6456] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6461:6456] * PIXEL_SIZE && v_count < i_worm_y[6461:6456] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1077 < i_size && h_count >= i_worm_x[6467:6462] * PIXEL_SIZE && h_count < i_worm_x[6467:6462] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6467:6462] * PIXEL_SIZE && v_count < i_worm_y[6467:6462] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1078 < i_size && h_count >= i_worm_x[6473:6468] * PIXEL_SIZE && h_count < i_worm_x[6473:6468] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6473:6468] * PIXEL_SIZE && v_count < i_worm_y[6473:6468] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1079 < i_size && h_count >= i_worm_x[6479:6474] * PIXEL_SIZE && h_count < i_worm_x[6479:6474] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6479:6474] * PIXEL_SIZE && v_count < i_worm_y[6479:6474] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1080 < i_size && h_count >= i_worm_x[6485:6480] * PIXEL_SIZE && h_count < i_worm_x[6485:6480] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6485:6480] * PIXEL_SIZE && v_count < i_worm_y[6485:6480] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1081 < i_size && h_count >= i_worm_x[6491:6486] * PIXEL_SIZE && h_count < i_worm_x[6491:6486] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6491:6486] * PIXEL_SIZE && v_count < i_worm_y[6491:6486] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1082 < i_size && h_count >= i_worm_x[6497:6492] * PIXEL_SIZE && h_count < i_worm_x[6497:6492] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6497:6492] * PIXEL_SIZE && v_count < i_worm_y[6497:6492] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1083 < i_size && h_count >= i_worm_x[6503:6498] * PIXEL_SIZE && h_count < i_worm_x[6503:6498] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6503:6498] * PIXEL_SIZE && v_count < i_worm_y[6503:6498] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1084 < i_size && h_count >= i_worm_x[6509:6504] * PIXEL_SIZE && h_count < i_worm_x[6509:6504] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6509:6504] * PIXEL_SIZE && v_count < i_worm_y[6509:6504] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1085 < i_size && h_count >= i_worm_x[6515:6510] * PIXEL_SIZE && h_count < i_worm_x[6515:6510] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6515:6510] * PIXEL_SIZE && v_count < i_worm_y[6515:6510] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1086 < i_size && h_count >= i_worm_x[6521:6516] * PIXEL_SIZE && h_count < i_worm_x[6521:6516] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6521:6516] * PIXEL_SIZE && v_count < i_worm_y[6521:6516] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1087 < i_size && h_count >= i_worm_x[6527:6522] * PIXEL_SIZE && h_count < i_worm_x[6527:6522] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6527:6522] * PIXEL_SIZE && v_count < i_worm_y[6527:6522] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1088 < i_size && h_count >= i_worm_x[6533:6528] * PIXEL_SIZE && h_count < i_worm_x[6533:6528] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6533:6528] * PIXEL_SIZE && v_count < i_worm_y[6533:6528] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1089 < i_size && h_count >= i_worm_x[6539:6534] * PIXEL_SIZE && h_count < i_worm_x[6539:6534] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6539:6534] * PIXEL_SIZE && v_count < i_worm_y[6539:6534] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1090 < i_size && h_count >= i_worm_x[6545:6540] * PIXEL_SIZE && h_count < i_worm_x[6545:6540] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6545:6540] * PIXEL_SIZE && v_count < i_worm_y[6545:6540] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1091 < i_size && h_count >= i_worm_x[6551:6546] * PIXEL_SIZE && h_count < i_worm_x[6551:6546] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6551:6546] * PIXEL_SIZE && v_count < i_worm_y[6551:6546] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1092 < i_size && h_count >= i_worm_x[6557:6552] * PIXEL_SIZE && h_count < i_worm_x[6557:6552] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6557:6552] * PIXEL_SIZE && v_count < i_worm_y[6557:6552] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1093 < i_size && h_count >= i_worm_x[6563:6558] * PIXEL_SIZE && h_count < i_worm_x[6563:6558] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6563:6558] * PIXEL_SIZE && v_count < i_worm_y[6563:6558] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1094 < i_size && h_count >= i_worm_x[6569:6564] * PIXEL_SIZE && h_count < i_worm_x[6569:6564] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6569:6564] * PIXEL_SIZE && v_count < i_worm_y[6569:6564] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1095 < i_size && h_count >= i_worm_x[6575:6570] * PIXEL_SIZE && h_count < i_worm_x[6575:6570] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6575:6570] * PIXEL_SIZE && v_count < i_worm_y[6575:6570] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1096 < i_size && h_count >= i_worm_x[6581:6576] * PIXEL_SIZE && h_count < i_worm_x[6581:6576] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6581:6576] * PIXEL_SIZE && v_count < i_worm_y[6581:6576] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1097 < i_size && h_count >= i_worm_x[6587:6582] * PIXEL_SIZE && h_count < i_worm_x[6587:6582] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6587:6582] * PIXEL_SIZE && v_count < i_worm_y[6587:6582] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1098 < i_size && h_count >= i_worm_x[6593:6588] * PIXEL_SIZE && h_count < i_worm_x[6593:6588] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6593:6588] * PIXEL_SIZE && v_count < i_worm_y[6593:6588] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1099 < i_size && h_count >= i_worm_x[6599:6594] * PIXEL_SIZE && h_count < i_worm_x[6599:6594] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6599:6594] * PIXEL_SIZE && v_count < i_worm_y[6599:6594] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1100 < i_size && h_count >= i_worm_x[6605:6600] * PIXEL_SIZE && h_count < i_worm_x[6605:6600] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6605:6600] * PIXEL_SIZE && v_count < i_worm_y[6605:6600] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1101 < i_size && h_count >= i_worm_x[6611:6606] * PIXEL_SIZE && h_count < i_worm_x[6611:6606] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6611:6606] * PIXEL_SIZE && v_count < i_worm_y[6611:6606] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1102 < i_size && h_count >= i_worm_x[6617:6612] * PIXEL_SIZE && h_count < i_worm_x[6617:6612] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6617:6612] * PIXEL_SIZE && v_count < i_worm_y[6617:6612] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1103 < i_size && h_count >= i_worm_x[6623:6618] * PIXEL_SIZE && h_count < i_worm_x[6623:6618] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6623:6618] * PIXEL_SIZE && v_count < i_worm_y[6623:6618] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1104 < i_size && h_count >= i_worm_x[6629:6624] * PIXEL_SIZE && h_count < i_worm_x[6629:6624] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6629:6624] * PIXEL_SIZE && v_count < i_worm_y[6629:6624] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1105 < i_size && h_count >= i_worm_x[6635:6630] * PIXEL_SIZE && h_count < i_worm_x[6635:6630] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6635:6630] * PIXEL_SIZE && v_count < i_worm_y[6635:6630] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1106 < i_size && h_count >= i_worm_x[6641:6636] * PIXEL_SIZE && h_count < i_worm_x[6641:6636] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6641:6636] * PIXEL_SIZE && v_count < i_worm_y[6641:6636] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1107 < i_size && h_count >= i_worm_x[6647:6642] * PIXEL_SIZE && h_count < i_worm_x[6647:6642] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6647:6642] * PIXEL_SIZE && v_count < i_worm_y[6647:6642] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1108 < i_size && h_count >= i_worm_x[6653:6648] * PIXEL_SIZE && h_count < i_worm_x[6653:6648] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6653:6648] * PIXEL_SIZE && v_count < i_worm_y[6653:6648] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1109 < i_size && h_count >= i_worm_x[6659:6654] * PIXEL_SIZE && h_count < i_worm_x[6659:6654] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6659:6654] * PIXEL_SIZE && v_count < i_worm_y[6659:6654] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1110 < i_size && h_count >= i_worm_x[6665:6660] * PIXEL_SIZE && h_count < i_worm_x[6665:6660] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6665:6660] * PIXEL_SIZE && v_count < i_worm_y[6665:6660] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1111 < i_size && h_count >= i_worm_x[6671:6666] * PIXEL_SIZE && h_count < i_worm_x[6671:6666] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6671:6666] * PIXEL_SIZE && v_count < i_worm_y[6671:6666] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1112 < i_size && h_count >= i_worm_x[6677:6672] * PIXEL_SIZE && h_count < i_worm_x[6677:6672] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6677:6672] * PIXEL_SIZE && v_count < i_worm_y[6677:6672] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1113 < i_size && h_count >= i_worm_x[6683:6678] * PIXEL_SIZE && h_count < i_worm_x[6683:6678] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6683:6678] * PIXEL_SIZE && v_count < i_worm_y[6683:6678] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1114 < i_size && h_count >= i_worm_x[6689:6684] * PIXEL_SIZE && h_count < i_worm_x[6689:6684] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6689:6684] * PIXEL_SIZE && v_count < i_worm_y[6689:6684] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1115 < i_size && h_count >= i_worm_x[6695:6690] * PIXEL_SIZE && h_count < i_worm_x[6695:6690] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6695:6690] * PIXEL_SIZE && v_count < i_worm_y[6695:6690] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1116 < i_size && h_count >= i_worm_x[6701:6696] * PIXEL_SIZE && h_count < i_worm_x[6701:6696] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6701:6696] * PIXEL_SIZE && v_count < i_worm_y[6701:6696] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1117 < i_size && h_count >= i_worm_x[6707:6702] * PIXEL_SIZE && h_count < i_worm_x[6707:6702] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6707:6702] * PIXEL_SIZE && v_count < i_worm_y[6707:6702] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1118 < i_size && h_count >= i_worm_x[6713:6708] * PIXEL_SIZE && h_count < i_worm_x[6713:6708] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6713:6708] * PIXEL_SIZE && v_count < i_worm_y[6713:6708] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1119 < i_size && h_count >= i_worm_x[6719:6714] * PIXEL_SIZE && h_count < i_worm_x[6719:6714] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6719:6714] * PIXEL_SIZE && v_count < i_worm_y[6719:6714] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1120 < i_size && h_count >= i_worm_x[6725:6720] * PIXEL_SIZE && h_count < i_worm_x[6725:6720] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6725:6720] * PIXEL_SIZE && v_count < i_worm_y[6725:6720] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1121 < i_size && h_count >= i_worm_x[6731:6726] * PIXEL_SIZE && h_count < i_worm_x[6731:6726] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6731:6726] * PIXEL_SIZE && v_count < i_worm_y[6731:6726] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1122 < i_size && h_count >= i_worm_x[6737:6732] * PIXEL_SIZE && h_count < i_worm_x[6737:6732] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6737:6732] * PIXEL_SIZE && v_count < i_worm_y[6737:6732] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1123 < i_size && h_count >= i_worm_x[6743:6738] * PIXEL_SIZE && h_count < i_worm_x[6743:6738] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6743:6738] * PIXEL_SIZE && v_count < i_worm_y[6743:6738] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1124 < i_size && h_count >= i_worm_x[6749:6744] * PIXEL_SIZE && h_count < i_worm_x[6749:6744] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6749:6744] * PIXEL_SIZE && v_count < i_worm_y[6749:6744] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1125 < i_size && h_count >= i_worm_x[6755:6750] * PIXEL_SIZE && h_count < i_worm_x[6755:6750] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6755:6750] * PIXEL_SIZE && v_count < i_worm_y[6755:6750] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1126 < i_size && h_count >= i_worm_x[6761:6756] * PIXEL_SIZE && h_count < i_worm_x[6761:6756] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6761:6756] * PIXEL_SIZE && v_count < i_worm_y[6761:6756] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1127 < i_size && h_count >= i_worm_x[6767:6762] * PIXEL_SIZE && h_count < i_worm_x[6767:6762] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6767:6762] * PIXEL_SIZE && v_count < i_worm_y[6767:6762] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1128 < i_size && h_count >= i_worm_x[6773:6768] * PIXEL_SIZE && h_count < i_worm_x[6773:6768] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6773:6768] * PIXEL_SIZE && v_count < i_worm_y[6773:6768] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1129 < i_size && h_count >= i_worm_x[6779:6774] * PIXEL_SIZE && h_count < i_worm_x[6779:6774] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6779:6774] * PIXEL_SIZE && v_count < i_worm_y[6779:6774] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1130 < i_size && h_count >= i_worm_x[6785:6780] * PIXEL_SIZE && h_count < i_worm_x[6785:6780] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6785:6780] * PIXEL_SIZE && v_count < i_worm_y[6785:6780] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1131 < i_size && h_count >= i_worm_x[6791:6786] * PIXEL_SIZE && h_count < i_worm_x[6791:6786] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6791:6786] * PIXEL_SIZE && v_count < i_worm_y[6791:6786] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1132 < i_size && h_count >= i_worm_x[6797:6792] * PIXEL_SIZE && h_count < i_worm_x[6797:6792] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6797:6792] * PIXEL_SIZE && v_count < i_worm_y[6797:6792] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1133 < i_size && h_count >= i_worm_x[6803:6798] * PIXEL_SIZE && h_count < i_worm_x[6803:6798] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6803:6798] * PIXEL_SIZE && v_count < i_worm_y[6803:6798] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1134 < i_size && h_count >= i_worm_x[6809:6804] * PIXEL_SIZE && h_count < i_worm_x[6809:6804] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6809:6804] * PIXEL_SIZE && v_count < i_worm_y[6809:6804] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1135 < i_size && h_count >= i_worm_x[6815:6810] * PIXEL_SIZE && h_count < i_worm_x[6815:6810] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6815:6810] * PIXEL_SIZE && v_count < i_worm_y[6815:6810] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1136 < i_size && h_count >= i_worm_x[6821:6816] * PIXEL_SIZE && h_count < i_worm_x[6821:6816] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6821:6816] * PIXEL_SIZE && v_count < i_worm_y[6821:6816] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1137 < i_size && h_count >= i_worm_x[6827:6822] * PIXEL_SIZE && h_count < i_worm_x[6827:6822] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6827:6822] * PIXEL_SIZE && v_count < i_worm_y[6827:6822] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1138 < i_size && h_count >= i_worm_x[6833:6828] * PIXEL_SIZE && h_count < i_worm_x[6833:6828] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6833:6828] * PIXEL_SIZE && v_count < i_worm_y[6833:6828] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1139 < i_size && h_count >= i_worm_x[6839:6834] * PIXEL_SIZE && h_count < i_worm_x[6839:6834] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6839:6834] * PIXEL_SIZE && v_count < i_worm_y[6839:6834] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1140 < i_size && h_count >= i_worm_x[6845:6840] * PIXEL_SIZE && h_count < i_worm_x[6845:6840] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6845:6840] * PIXEL_SIZE && v_count < i_worm_y[6845:6840] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1141 < i_size && h_count >= i_worm_x[6851:6846] * PIXEL_SIZE && h_count < i_worm_x[6851:6846] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6851:6846] * PIXEL_SIZE && v_count < i_worm_y[6851:6846] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1142 < i_size && h_count >= i_worm_x[6857:6852] * PIXEL_SIZE && h_count < i_worm_x[6857:6852] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6857:6852] * PIXEL_SIZE && v_count < i_worm_y[6857:6852] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1143 < i_size && h_count >= i_worm_x[6863:6858] * PIXEL_SIZE && h_count < i_worm_x[6863:6858] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6863:6858] * PIXEL_SIZE && v_count < i_worm_y[6863:6858] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1144 < i_size && h_count >= i_worm_x[6869:6864] * PIXEL_SIZE && h_count < i_worm_x[6869:6864] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6869:6864] * PIXEL_SIZE && v_count < i_worm_y[6869:6864] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1145 < i_size && h_count >= i_worm_x[6875:6870] * PIXEL_SIZE && h_count < i_worm_x[6875:6870] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6875:6870] * PIXEL_SIZE && v_count < i_worm_y[6875:6870] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1146 < i_size && h_count >= i_worm_x[6881:6876] * PIXEL_SIZE && h_count < i_worm_x[6881:6876] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6881:6876] * PIXEL_SIZE && v_count < i_worm_y[6881:6876] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1147 < i_size && h_count >= i_worm_x[6887:6882] * PIXEL_SIZE && h_count < i_worm_x[6887:6882] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6887:6882] * PIXEL_SIZE && v_count < i_worm_y[6887:6882] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1148 < i_size && h_count >= i_worm_x[6893:6888] * PIXEL_SIZE && h_count < i_worm_x[6893:6888] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6893:6888] * PIXEL_SIZE && v_count < i_worm_y[6893:6888] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1149 < i_size && h_count >= i_worm_x[6899:6894] * PIXEL_SIZE && h_count < i_worm_x[6899:6894] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6899:6894] * PIXEL_SIZE && v_count < i_worm_y[6899:6894] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1150 < i_size && h_count >= i_worm_x[6905:6900] * PIXEL_SIZE && h_count < i_worm_x[6905:6900] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6905:6900] * PIXEL_SIZE && v_count < i_worm_y[6905:6900] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1151 < i_size && h_count >= i_worm_x[6911:6906] * PIXEL_SIZE && h_count < i_worm_x[6911:6906] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6911:6906] * PIXEL_SIZE && v_count < i_worm_y[6911:6906] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1152 < i_size && h_count >= i_worm_x[6917:6912] * PIXEL_SIZE && h_count < i_worm_x[6917:6912] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6917:6912] * PIXEL_SIZE && v_count < i_worm_y[6917:6912] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1153 < i_size && h_count >= i_worm_x[6923:6918] * PIXEL_SIZE && h_count < i_worm_x[6923:6918] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6923:6918] * PIXEL_SIZE && v_count < i_worm_y[6923:6918] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1154 < i_size && h_count >= i_worm_x[6929:6924] * PIXEL_SIZE && h_count < i_worm_x[6929:6924] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6929:6924] * PIXEL_SIZE && v_count < i_worm_y[6929:6924] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1155 < i_size && h_count >= i_worm_x[6935:6930] * PIXEL_SIZE && h_count < i_worm_x[6935:6930] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6935:6930] * PIXEL_SIZE && v_count < i_worm_y[6935:6930] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1156 < i_size && h_count >= i_worm_x[6941:6936] * PIXEL_SIZE && h_count < i_worm_x[6941:6936] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6941:6936] * PIXEL_SIZE && v_count < i_worm_y[6941:6936] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1157 < i_size && h_count >= i_worm_x[6947:6942] * PIXEL_SIZE && h_count < i_worm_x[6947:6942] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6947:6942] * PIXEL_SIZE && v_count < i_worm_y[6947:6942] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1158 < i_size && h_count >= i_worm_x[6953:6948] * PIXEL_SIZE && h_count < i_worm_x[6953:6948] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6953:6948] * PIXEL_SIZE && v_count < i_worm_y[6953:6948] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1159 < i_size && h_count >= i_worm_x[6959:6954] * PIXEL_SIZE && h_count < i_worm_x[6959:6954] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6959:6954] * PIXEL_SIZE && v_count < i_worm_y[6959:6954] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1160 < i_size && h_count >= i_worm_x[6965:6960] * PIXEL_SIZE && h_count < i_worm_x[6965:6960] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6965:6960] * PIXEL_SIZE && v_count < i_worm_y[6965:6960] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1161 < i_size && h_count >= i_worm_x[6971:6966] * PIXEL_SIZE && h_count < i_worm_x[6971:6966] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6971:6966] * PIXEL_SIZE && v_count < i_worm_y[6971:6966] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1162 < i_size && h_count >= i_worm_x[6977:6972] * PIXEL_SIZE && h_count < i_worm_x[6977:6972] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6977:6972] * PIXEL_SIZE && v_count < i_worm_y[6977:6972] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1163 < i_size && h_count >= i_worm_x[6983:6978] * PIXEL_SIZE && h_count < i_worm_x[6983:6978] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6983:6978] * PIXEL_SIZE && v_count < i_worm_y[6983:6978] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1164 < i_size && h_count >= i_worm_x[6989:6984] * PIXEL_SIZE && h_count < i_worm_x[6989:6984] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6989:6984] * PIXEL_SIZE && v_count < i_worm_y[6989:6984] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1165 < i_size && h_count >= i_worm_x[6995:6990] * PIXEL_SIZE && h_count < i_worm_x[6995:6990] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[6995:6990] * PIXEL_SIZE && v_count < i_worm_y[6995:6990] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1166 < i_size && h_count >= i_worm_x[7001:6996] * PIXEL_SIZE && h_count < i_worm_x[7001:6996] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7001:6996] * PIXEL_SIZE && v_count < i_worm_y[7001:6996] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1167 < i_size && h_count >= i_worm_x[7007:7002] * PIXEL_SIZE && h_count < i_worm_x[7007:7002] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7007:7002] * PIXEL_SIZE && v_count < i_worm_y[7007:7002] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1168 < i_size && h_count >= i_worm_x[7013:7008] * PIXEL_SIZE && h_count < i_worm_x[7013:7008] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7013:7008] * PIXEL_SIZE && v_count < i_worm_y[7013:7008] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1169 < i_size && h_count >= i_worm_x[7019:7014] * PIXEL_SIZE && h_count < i_worm_x[7019:7014] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7019:7014] * PIXEL_SIZE && v_count < i_worm_y[7019:7014] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1170 < i_size && h_count >= i_worm_x[7025:7020] * PIXEL_SIZE && h_count < i_worm_x[7025:7020] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7025:7020] * PIXEL_SIZE && v_count < i_worm_y[7025:7020] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1171 < i_size && h_count >= i_worm_x[7031:7026] * PIXEL_SIZE && h_count < i_worm_x[7031:7026] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7031:7026] * PIXEL_SIZE && v_count < i_worm_y[7031:7026] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1172 < i_size && h_count >= i_worm_x[7037:7032] * PIXEL_SIZE && h_count < i_worm_x[7037:7032] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7037:7032] * PIXEL_SIZE && v_count < i_worm_y[7037:7032] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1173 < i_size && h_count >= i_worm_x[7043:7038] * PIXEL_SIZE && h_count < i_worm_x[7043:7038] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7043:7038] * PIXEL_SIZE && v_count < i_worm_y[7043:7038] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1174 < i_size && h_count >= i_worm_x[7049:7044] * PIXEL_SIZE && h_count < i_worm_x[7049:7044] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7049:7044] * PIXEL_SIZE && v_count < i_worm_y[7049:7044] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1175 < i_size && h_count >= i_worm_x[7055:7050] * PIXEL_SIZE && h_count < i_worm_x[7055:7050] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7055:7050] * PIXEL_SIZE && v_count < i_worm_y[7055:7050] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1176 < i_size && h_count >= i_worm_x[7061:7056] * PIXEL_SIZE && h_count < i_worm_x[7061:7056] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7061:7056] * PIXEL_SIZE && v_count < i_worm_y[7061:7056] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1177 < i_size && h_count >= i_worm_x[7067:7062] * PIXEL_SIZE && h_count < i_worm_x[7067:7062] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7067:7062] * PIXEL_SIZE && v_count < i_worm_y[7067:7062] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1178 < i_size && h_count >= i_worm_x[7073:7068] * PIXEL_SIZE && h_count < i_worm_x[7073:7068] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7073:7068] * PIXEL_SIZE && v_count < i_worm_y[7073:7068] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1179 < i_size && h_count >= i_worm_x[7079:7074] * PIXEL_SIZE && h_count < i_worm_x[7079:7074] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7079:7074] * PIXEL_SIZE && v_count < i_worm_y[7079:7074] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1180 < i_size && h_count >= i_worm_x[7085:7080] * PIXEL_SIZE && h_count < i_worm_x[7085:7080] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7085:7080] * PIXEL_SIZE && v_count < i_worm_y[7085:7080] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1181 < i_size && h_count >= i_worm_x[7091:7086] * PIXEL_SIZE && h_count < i_worm_x[7091:7086] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7091:7086] * PIXEL_SIZE && v_count < i_worm_y[7091:7086] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1182 < i_size && h_count >= i_worm_x[7097:7092] * PIXEL_SIZE && h_count < i_worm_x[7097:7092] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7097:7092] * PIXEL_SIZE && v_count < i_worm_y[7097:7092] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1183 < i_size && h_count >= i_worm_x[7103:7098] * PIXEL_SIZE && h_count < i_worm_x[7103:7098] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7103:7098] * PIXEL_SIZE && v_count < i_worm_y[7103:7098] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1184 < i_size && h_count >= i_worm_x[7109:7104] * PIXEL_SIZE && h_count < i_worm_x[7109:7104] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7109:7104] * PIXEL_SIZE && v_count < i_worm_y[7109:7104] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1185 < i_size && h_count >= i_worm_x[7115:7110] * PIXEL_SIZE && h_count < i_worm_x[7115:7110] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7115:7110] * PIXEL_SIZE && v_count < i_worm_y[7115:7110] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1186 < i_size && h_count >= i_worm_x[7121:7116] * PIXEL_SIZE && h_count < i_worm_x[7121:7116] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7121:7116] * PIXEL_SIZE && v_count < i_worm_y[7121:7116] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1187 < i_size && h_count >= i_worm_x[7127:7122] * PIXEL_SIZE && h_count < i_worm_x[7127:7122] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7127:7122] * PIXEL_SIZE && v_count < i_worm_y[7127:7122] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1188 < i_size && h_count >= i_worm_x[7133:7128] * PIXEL_SIZE && h_count < i_worm_x[7133:7128] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7133:7128] * PIXEL_SIZE && v_count < i_worm_y[7133:7128] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1189 < i_size && h_count >= i_worm_x[7139:7134] * PIXEL_SIZE && h_count < i_worm_x[7139:7134] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7139:7134] * PIXEL_SIZE && v_count < i_worm_y[7139:7134] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1190 < i_size && h_count >= i_worm_x[7145:7140] * PIXEL_SIZE && h_count < i_worm_x[7145:7140] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7145:7140] * PIXEL_SIZE && v_count < i_worm_y[7145:7140] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1191 < i_size && h_count >= i_worm_x[7151:7146] * PIXEL_SIZE && h_count < i_worm_x[7151:7146] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7151:7146] * PIXEL_SIZE && v_count < i_worm_y[7151:7146] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1192 < i_size && h_count >= i_worm_x[7157:7152] * PIXEL_SIZE && h_count < i_worm_x[7157:7152] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7157:7152] * PIXEL_SIZE && v_count < i_worm_y[7157:7152] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1193 < i_size && h_count >= i_worm_x[7163:7158] * PIXEL_SIZE && h_count < i_worm_x[7163:7158] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7163:7158] * PIXEL_SIZE && v_count < i_worm_y[7163:7158] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1194 < i_size && h_count >= i_worm_x[7169:7164] * PIXEL_SIZE && h_count < i_worm_x[7169:7164] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7169:7164] * PIXEL_SIZE && v_count < i_worm_y[7169:7164] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1195 < i_size && h_count >= i_worm_x[7175:7170] * PIXEL_SIZE && h_count < i_worm_x[7175:7170] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7175:7170] * PIXEL_SIZE && v_count < i_worm_y[7175:7170] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1196 < i_size && h_count >= i_worm_x[7181:7176] * PIXEL_SIZE && h_count < i_worm_x[7181:7176] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7181:7176] * PIXEL_SIZE && v_count < i_worm_y[7181:7176] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1197 < i_size && h_count >= i_worm_x[7187:7182] * PIXEL_SIZE && h_count < i_worm_x[7187:7182] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7187:7182] * PIXEL_SIZE && v_count < i_worm_y[7187:7182] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1198 < i_size && h_count >= i_worm_x[7193:7188] * PIXEL_SIZE && h_count < i_worm_x[7193:7188] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7193:7188] * PIXEL_SIZE && v_count < i_worm_y[7193:7188] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1199 < i_size && h_count >= i_worm_x[7199:7194] * PIXEL_SIZE && h_count < i_worm_x[7199:7194] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7199:7194] * PIXEL_SIZE && v_count < i_worm_y[7199:7194] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1200 < i_size && h_count >= i_worm_x[7205:7200] * PIXEL_SIZE && h_count < i_worm_x[7205:7200] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7205:7200] * PIXEL_SIZE && v_count < i_worm_y[7205:7200] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1201 < i_size && h_count >= i_worm_x[7211:7206] * PIXEL_SIZE && h_count < i_worm_x[7211:7206] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7211:7206] * PIXEL_SIZE && v_count < i_worm_y[7211:7206] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1202 < i_size && h_count >= i_worm_x[7217:7212] * PIXEL_SIZE && h_count < i_worm_x[7217:7212] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7217:7212] * PIXEL_SIZE && v_count < i_worm_y[7217:7212] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1203 < i_size && h_count >= i_worm_x[7223:7218] * PIXEL_SIZE && h_count < i_worm_x[7223:7218] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7223:7218] * PIXEL_SIZE && v_count < i_worm_y[7223:7218] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1204 < i_size && h_count >= i_worm_x[7229:7224] * PIXEL_SIZE && h_count < i_worm_x[7229:7224] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7229:7224] * PIXEL_SIZE && v_count < i_worm_y[7229:7224] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1205 < i_size && h_count >= i_worm_x[7235:7230] * PIXEL_SIZE && h_count < i_worm_x[7235:7230] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7235:7230] * PIXEL_SIZE && v_count < i_worm_y[7235:7230] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1206 < i_size && h_count >= i_worm_x[7241:7236] * PIXEL_SIZE && h_count < i_worm_x[7241:7236] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7241:7236] * PIXEL_SIZE && v_count < i_worm_y[7241:7236] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1207 < i_size && h_count >= i_worm_x[7247:7242] * PIXEL_SIZE && h_count < i_worm_x[7247:7242] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7247:7242] * PIXEL_SIZE && v_count < i_worm_y[7247:7242] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1208 < i_size && h_count >= i_worm_x[7253:7248] * PIXEL_SIZE && h_count < i_worm_x[7253:7248] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7253:7248] * PIXEL_SIZE && v_count < i_worm_y[7253:7248] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1209 < i_size && h_count >= i_worm_x[7259:7254] * PIXEL_SIZE && h_count < i_worm_x[7259:7254] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7259:7254] * PIXEL_SIZE && v_count < i_worm_y[7259:7254] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1210 < i_size && h_count >= i_worm_x[7265:7260] * PIXEL_SIZE && h_count < i_worm_x[7265:7260] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7265:7260] * PIXEL_SIZE && v_count < i_worm_y[7265:7260] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1211 < i_size && h_count >= i_worm_x[7271:7266] * PIXEL_SIZE && h_count < i_worm_x[7271:7266] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7271:7266] * PIXEL_SIZE && v_count < i_worm_y[7271:7266] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1212 < i_size && h_count >= i_worm_x[7277:7272] * PIXEL_SIZE && h_count < i_worm_x[7277:7272] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7277:7272] * PIXEL_SIZE && v_count < i_worm_y[7277:7272] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1213 < i_size && h_count >= i_worm_x[7283:7278] * PIXEL_SIZE && h_count < i_worm_x[7283:7278] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7283:7278] * PIXEL_SIZE && v_count < i_worm_y[7283:7278] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1214 < i_size && h_count >= i_worm_x[7289:7284] * PIXEL_SIZE && h_count < i_worm_x[7289:7284] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7289:7284] * PIXEL_SIZE && v_count < i_worm_y[7289:7284] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1215 < i_size && h_count >= i_worm_x[7295:7290] * PIXEL_SIZE && h_count < i_worm_x[7295:7290] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7295:7290] * PIXEL_SIZE && v_count < i_worm_y[7295:7290] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1216 < i_size && h_count >= i_worm_x[7301:7296] * PIXEL_SIZE && h_count < i_worm_x[7301:7296] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7301:7296] * PIXEL_SIZE && v_count < i_worm_y[7301:7296] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1217 < i_size && h_count >= i_worm_x[7307:7302] * PIXEL_SIZE && h_count < i_worm_x[7307:7302] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7307:7302] * PIXEL_SIZE && v_count < i_worm_y[7307:7302] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1218 < i_size && h_count >= i_worm_x[7313:7308] * PIXEL_SIZE && h_count < i_worm_x[7313:7308] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7313:7308] * PIXEL_SIZE && v_count < i_worm_y[7313:7308] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1219 < i_size && h_count >= i_worm_x[7319:7314] * PIXEL_SIZE && h_count < i_worm_x[7319:7314] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7319:7314] * PIXEL_SIZE && v_count < i_worm_y[7319:7314] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1220 < i_size && h_count >= i_worm_x[7325:7320] * PIXEL_SIZE && h_count < i_worm_x[7325:7320] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7325:7320] * PIXEL_SIZE && v_count < i_worm_y[7325:7320] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1221 < i_size && h_count >= i_worm_x[7331:7326] * PIXEL_SIZE && h_count < i_worm_x[7331:7326] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7331:7326] * PIXEL_SIZE && v_count < i_worm_y[7331:7326] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1222 < i_size && h_count >= i_worm_x[7337:7332] * PIXEL_SIZE && h_count < i_worm_x[7337:7332] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7337:7332] * PIXEL_SIZE && v_count < i_worm_y[7337:7332] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1223 < i_size && h_count >= i_worm_x[7343:7338] * PIXEL_SIZE && h_count < i_worm_x[7343:7338] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7343:7338] * PIXEL_SIZE && v_count < i_worm_y[7343:7338] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1224 < i_size && h_count >= i_worm_x[7349:7344] * PIXEL_SIZE && h_count < i_worm_x[7349:7344] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7349:7344] * PIXEL_SIZE && v_count < i_worm_y[7349:7344] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1225 < i_size && h_count >= i_worm_x[7355:7350] * PIXEL_SIZE && h_count < i_worm_x[7355:7350] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7355:7350] * PIXEL_SIZE && v_count < i_worm_y[7355:7350] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1226 < i_size && h_count >= i_worm_x[7361:7356] * PIXEL_SIZE && h_count < i_worm_x[7361:7356] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7361:7356] * PIXEL_SIZE && v_count < i_worm_y[7361:7356] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1227 < i_size && h_count >= i_worm_x[7367:7362] * PIXEL_SIZE && h_count < i_worm_x[7367:7362] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7367:7362] * PIXEL_SIZE && v_count < i_worm_y[7367:7362] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1228 < i_size && h_count >= i_worm_x[7373:7368] * PIXEL_SIZE && h_count < i_worm_x[7373:7368] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7373:7368] * PIXEL_SIZE && v_count < i_worm_y[7373:7368] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1229 < i_size && h_count >= i_worm_x[7379:7374] * PIXEL_SIZE && h_count < i_worm_x[7379:7374] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7379:7374] * PIXEL_SIZE && v_count < i_worm_y[7379:7374] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1230 < i_size && h_count >= i_worm_x[7385:7380] * PIXEL_SIZE && h_count < i_worm_x[7385:7380] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7385:7380] * PIXEL_SIZE && v_count < i_worm_y[7385:7380] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1231 < i_size && h_count >= i_worm_x[7391:7386] * PIXEL_SIZE && h_count < i_worm_x[7391:7386] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7391:7386] * PIXEL_SIZE && v_count < i_worm_y[7391:7386] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1232 < i_size && h_count >= i_worm_x[7397:7392] * PIXEL_SIZE && h_count < i_worm_x[7397:7392] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7397:7392] * PIXEL_SIZE && v_count < i_worm_y[7397:7392] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1233 < i_size && h_count >= i_worm_x[7403:7398] * PIXEL_SIZE && h_count < i_worm_x[7403:7398] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7403:7398] * PIXEL_SIZE && v_count < i_worm_y[7403:7398] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1234 < i_size && h_count >= i_worm_x[7409:7404] * PIXEL_SIZE && h_count < i_worm_x[7409:7404] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7409:7404] * PIXEL_SIZE && v_count < i_worm_y[7409:7404] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1235 < i_size && h_count >= i_worm_x[7415:7410] * PIXEL_SIZE && h_count < i_worm_x[7415:7410] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7415:7410] * PIXEL_SIZE && v_count < i_worm_y[7415:7410] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1236 < i_size && h_count >= i_worm_x[7421:7416] * PIXEL_SIZE && h_count < i_worm_x[7421:7416] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7421:7416] * PIXEL_SIZE && v_count < i_worm_y[7421:7416] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1237 < i_size && h_count >= i_worm_x[7427:7422] * PIXEL_SIZE && h_count < i_worm_x[7427:7422] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7427:7422] * PIXEL_SIZE && v_count < i_worm_y[7427:7422] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1238 < i_size && h_count >= i_worm_x[7433:7428] * PIXEL_SIZE && h_count < i_worm_x[7433:7428] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7433:7428] * PIXEL_SIZE && v_count < i_worm_y[7433:7428] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1239 < i_size && h_count >= i_worm_x[7439:7434] * PIXEL_SIZE && h_count < i_worm_x[7439:7434] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7439:7434] * PIXEL_SIZE && v_count < i_worm_y[7439:7434] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1240 < i_size && h_count >= i_worm_x[7445:7440] * PIXEL_SIZE && h_count < i_worm_x[7445:7440] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7445:7440] * PIXEL_SIZE && v_count < i_worm_y[7445:7440] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1241 < i_size && h_count >= i_worm_x[7451:7446] * PIXEL_SIZE && h_count < i_worm_x[7451:7446] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7451:7446] * PIXEL_SIZE && v_count < i_worm_y[7451:7446] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1242 < i_size && h_count >= i_worm_x[7457:7452] * PIXEL_SIZE && h_count < i_worm_x[7457:7452] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7457:7452] * PIXEL_SIZE && v_count < i_worm_y[7457:7452] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1243 < i_size && h_count >= i_worm_x[7463:7458] * PIXEL_SIZE && h_count < i_worm_x[7463:7458] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7463:7458] * PIXEL_SIZE && v_count < i_worm_y[7463:7458] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1244 < i_size && h_count >= i_worm_x[7469:7464] * PIXEL_SIZE && h_count < i_worm_x[7469:7464] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7469:7464] * PIXEL_SIZE && v_count < i_worm_y[7469:7464] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1245 < i_size && h_count >= i_worm_x[7475:7470] * PIXEL_SIZE && h_count < i_worm_x[7475:7470] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7475:7470] * PIXEL_SIZE && v_count < i_worm_y[7475:7470] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1246 < i_size && h_count >= i_worm_x[7481:7476] * PIXEL_SIZE && h_count < i_worm_x[7481:7476] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7481:7476] * PIXEL_SIZE && v_count < i_worm_y[7481:7476] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1247 < i_size && h_count >= i_worm_x[7487:7482] * PIXEL_SIZE && h_count < i_worm_x[7487:7482] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7487:7482] * PIXEL_SIZE && v_count < i_worm_y[7487:7482] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1248 < i_size && h_count >= i_worm_x[7493:7488] * PIXEL_SIZE && h_count < i_worm_x[7493:7488] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7493:7488] * PIXEL_SIZE && v_count < i_worm_y[7493:7488] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1249 < i_size && h_count >= i_worm_x[7499:7494] * PIXEL_SIZE && h_count < i_worm_x[7499:7494] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7499:7494] * PIXEL_SIZE && v_count < i_worm_y[7499:7494] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1250 < i_size && h_count >= i_worm_x[7505:7500] * PIXEL_SIZE && h_count < i_worm_x[7505:7500] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7505:7500] * PIXEL_SIZE && v_count < i_worm_y[7505:7500] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1251 < i_size && h_count >= i_worm_x[7511:7506] * PIXEL_SIZE && h_count < i_worm_x[7511:7506] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7511:7506] * PIXEL_SIZE && v_count < i_worm_y[7511:7506] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1252 < i_size && h_count >= i_worm_x[7517:7512] * PIXEL_SIZE && h_count < i_worm_x[7517:7512] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7517:7512] * PIXEL_SIZE && v_count < i_worm_y[7517:7512] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1253 < i_size && h_count >= i_worm_x[7523:7518] * PIXEL_SIZE && h_count < i_worm_x[7523:7518] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7523:7518] * PIXEL_SIZE && v_count < i_worm_y[7523:7518] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1254 < i_size && h_count >= i_worm_x[7529:7524] * PIXEL_SIZE && h_count < i_worm_x[7529:7524] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7529:7524] * PIXEL_SIZE && v_count < i_worm_y[7529:7524] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1255 < i_size && h_count >= i_worm_x[7535:7530] * PIXEL_SIZE && h_count < i_worm_x[7535:7530] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7535:7530] * PIXEL_SIZE && v_count < i_worm_y[7535:7530] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1256 < i_size && h_count >= i_worm_x[7541:7536] * PIXEL_SIZE && h_count < i_worm_x[7541:7536] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7541:7536] * PIXEL_SIZE && v_count < i_worm_y[7541:7536] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1257 < i_size && h_count >= i_worm_x[7547:7542] * PIXEL_SIZE && h_count < i_worm_x[7547:7542] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7547:7542] * PIXEL_SIZE && v_count < i_worm_y[7547:7542] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1258 < i_size && h_count >= i_worm_x[7553:7548] * PIXEL_SIZE && h_count < i_worm_x[7553:7548] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7553:7548] * PIXEL_SIZE && v_count < i_worm_y[7553:7548] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1259 < i_size && h_count >= i_worm_x[7559:7554] * PIXEL_SIZE && h_count < i_worm_x[7559:7554] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7559:7554] * PIXEL_SIZE && v_count < i_worm_y[7559:7554] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1260 < i_size && h_count >= i_worm_x[7565:7560] * PIXEL_SIZE && h_count < i_worm_x[7565:7560] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7565:7560] * PIXEL_SIZE && v_count < i_worm_y[7565:7560] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1261 < i_size && h_count >= i_worm_x[7571:7566] * PIXEL_SIZE && h_count < i_worm_x[7571:7566] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7571:7566] * PIXEL_SIZE && v_count < i_worm_y[7571:7566] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1262 < i_size && h_count >= i_worm_x[7577:7572] * PIXEL_SIZE && h_count < i_worm_x[7577:7572] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7577:7572] * PIXEL_SIZE && v_count < i_worm_y[7577:7572] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1263 < i_size && h_count >= i_worm_x[7583:7578] * PIXEL_SIZE && h_count < i_worm_x[7583:7578] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7583:7578] * PIXEL_SIZE && v_count < i_worm_y[7583:7578] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1264 < i_size && h_count >= i_worm_x[7589:7584] * PIXEL_SIZE && h_count < i_worm_x[7589:7584] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7589:7584] * PIXEL_SIZE && v_count < i_worm_y[7589:7584] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1265 < i_size && h_count >= i_worm_x[7595:7590] * PIXEL_SIZE && h_count < i_worm_x[7595:7590] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7595:7590] * PIXEL_SIZE && v_count < i_worm_y[7595:7590] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1266 < i_size && h_count >= i_worm_x[7601:7596] * PIXEL_SIZE && h_count < i_worm_x[7601:7596] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7601:7596] * PIXEL_SIZE && v_count < i_worm_y[7601:7596] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1267 < i_size && h_count >= i_worm_x[7607:7602] * PIXEL_SIZE && h_count < i_worm_x[7607:7602] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7607:7602] * PIXEL_SIZE && v_count < i_worm_y[7607:7602] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1268 < i_size && h_count >= i_worm_x[7613:7608] * PIXEL_SIZE && h_count < i_worm_x[7613:7608] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7613:7608] * PIXEL_SIZE && v_count < i_worm_y[7613:7608] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1269 < i_size && h_count >= i_worm_x[7619:7614] * PIXEL_SIZE && h_count < i_worm_x[7619:7614] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7619:7614] * PIXEL_SIZE && v_count < i_worm_y[7619:7614] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1270 < i_size && h_count >= i_worm_x[7625:7620] * PIXEL_SIZE && h_count < i_worm_x[7625:7620] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7625:7620] * PIXEL_SIZE && v_count < i_worm_y[7625:7620] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1271 < i_size && h_count >= i_worm_x[7631:7626] * PIXEL_SIZE && h_count < i_worm_x[7631:7626] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7631:7626] * PIXEL_SIZE && v_count < i_worm_y[7631:7626] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1272 < i_size && h_count >= i_worm_x[7637:7632] * PIXEL_SIZE && h_count < i_worm_x[7637:7632] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7637:7632] * PIXEL_SIZE && v_count < i_worm_y[7637:7632] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1273 < i_size && h_count >= i_worm_x[7643:7638] * PIXEL_SIZE && h_count < i_worm_x[7643:7638] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7643:7638] * PIXEL_SIZE && v_count < i_worm_y[7643:7638] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1274 < i_size && h_count >= i_worm_x[7649:7644] * PIXEL_SIZE && h_count < i_worm_x[7649:7644] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7649:7644] * PIXEL_SIZE && v_count < i_worm_y[7649:7644] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1275 < i_size && h_count >= i_worm_x[7655:7650] * PIXEL_SIZE && h_count < i_worm_x[7655:7650] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7655:7650] * PIXEL_SIZE && v_count < i_worm_y[7655:7650] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1276 < i_size && h_count >= i_worm_x[7661:7656] * PIXEL_SIZE && h_count < i_worm_x[7661:7656] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7661:7656] * PIXEL_SIZE && v_count < i_worm_y[7661:7656] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1277 < i_size && h_count >= i_worm_x[7667:7662] * PIXEL_SIZE && h_count < i_worm_x[7667:7662] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7667:7662] * PIXEL_SIZE && v_count < i_worm_y[7667:7662] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1278 < i_size && h_count >= i_worm_x[7673:7668] * PIXEL_SIZE && h_count < i_worm_x[7673:7668] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7673:7668] * PIXEL_SIZE && v_count < i_worm_y[7673:7668] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1279 < i_size && h_count >= i_worm_x[7679:7674] * PIXEL_SIZE && h_count < i_worm_x[7679:7674] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7679:7674] * PIXEL_SIZE && v_count < i_worm_y[7679:7674] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1280 < i_size && h_count >= i_worm_x[7685:7680] * PIXEL_SIZE && h_count < i_worm_x[7685:7680] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7685:7680] * PIXEL_SIZE && v_count < i_worm_y[7685:7680] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1281 < i_size && h_count >= i_worm_x[7691:7686] * PIXEL_SIZE && h_count < i_worm_x[7691:7686] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7691:7686] * PIXEL_SIZE && v_count < i_worm_y[7691:7686] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1282 < i_size && h_count >= i_worm_x[7697:7692] * PIXEL_SIZE && h_count < i_worm_x[7697:7692] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7697:7692] * PIXEL_SIZE && v_count < i_worm_y[7697:7692] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1283 < i_size && h_count >= i_worm_x[7703:7698] * PIXEL_SIZE && h_count < i_worm_x[7703:7698] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7703:7698] * PIXEL_SIZE && v_count < i_worm_y[7703:7698] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1284 < i_size && h_count >= i_worm_x[7709:7704] * PIXEL_SIZE && h_count < i_worm_x[7709:7704] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7709:7704] * PIXEL_SIZE && v_count < i_worm_y[7709:7704] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1285 < i_size && h_count >= i_worm_x[7715:7710] * PIXEL_SIZE && h_count < i_worm_x[7715:7710] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7715:7710] * PIXEL_SIZE && v_count < i_worm_y[7715:7710] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1286 < i_size && h_count >= i_worm_x[7721:7716] * PIXEL_SIZE && h_count < i_worm_x[7721:7716] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7721:7716] * PIXEL_SIZE && v_count < i_worm_y[7721:7716] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1287 < i_size && h_count >= i_worm_x[7727:7722] * PIXEL_SIZE && h_count < i_worm_x[7727:7722] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7727:7722] * PIXEL_SIZE && v_count < i_worm_y[7727:7722] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1288 < i_size && h_count >= i_worm_x[7733:7728] * PIXEL_SIZE && h_count < i_worm_x[7733:7728] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7733:7728] * PIXEL_SIZE && v_count < i_worm_y[7733:7728] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1289 < i_size && h_count >= i_worm_x[7739:7734] * PIXEL_SIZE && h_count < i_worm_x[7739:7734] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7739:7734] * PIXEL_SIZE && v_count < i_worm_y[7739:7734] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1290 < i_size && h_count >= i_worm_x[7745:7740] * PIXEL_SIZE && h_count < i_worm_x[7745:7740] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7745:7740] * PIXEL_SIZE && v_count < i_worm_y[7745:7740] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1291 < i_size && h_count >= i_worm_x[7751:7746] * PIXEL_SIZE && h_count < i_worm_x[7751:7746] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7751:7746] * PIXEL_SIZE && v_count < i_worm_y[7751:7746] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1292 < i_size && h_count >= i_worm_x[7757:7752] * PIXEL_SIZE && h_count < i_worm_x[7757:7752] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7757:7752] * PIXEL_SIZE && v_count < i_worm_y[7757:7752] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1293 < i_size && h_count >= i_worm_x[7763:7758] * PIXEL_SIZE && h_count < i_worm_x[7763:7758] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7763:7758] * PIXEL_SIZE && v_count < i_worm_y[7763:7758] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1294 < i_size && h_count >= i_worm_x[7769:7764] * PIXEL_SIZE && h_count < i_worm_x[7769:7764] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7769:7764] * PIXEL_SIZE && v_count < i_worm_y[7769:7764] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1295 < i_size && h_count >= i_worm_x[7775:7770] * PIXEL_SIZE && h_count < i_worm_x[7775:7770] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7775:7770] * PIXEL_SIZE && v_count < i_worm_y[7775:7770] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1296 < i_size && h_count >= i_worm_x[7781:7776] * PIXEL_SIZE && h_count < i_worm_x[7781:7776] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7781:7776] * PIXEL_SIZE && v_count < i_worm_y[7781:7776] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1297 < i_size && h_count >= i_worm_x[7787:7782] * PIXEL_SIZE && h_count < i_worm_x[7787:7782] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7787:7782] * PIXEL_SIZE && v_count < i_worm_y[7787:7782] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1298 < i_size && h_count >= i_worm_x[7793:7788] * PIXEL_SIZE && h_count < i_worm_x[7793:7788] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7793:7788] * PIXEL_SIZE && v_count < i_worm_y[7793:7788] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1299 < i_size && h_count >= i_worm_x[7799:7794] * PIXEL_SIZE && h_count < i_worm_x[7799:7794] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7799:7794] * PIXEL_SIZE && v_count < i_worm_y[7799:7794] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1300 < i_size && h_count >= i_worm_x[7805:7800] * PIXEL_SIZE && h_count < i_worm_x[7805:7800] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7805:7800] * PIXEL_SIZE && v_count < i_worm_y[7805:7800] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1301 < i_size && h_count >= i_worm_x[7811:7806] * PIXEL_SIZE && h_count < i_worm_x[7811:7806] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7811:7806] * PIXEL_SIZE && v_count < i_worm_y[7811:7806] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1302 < i_size && h_count >= i_worm_x[7817:7812] * PIXEL_SIZE && h_count < i_worm_x[7817:7812] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7817:7812] * PIXEL_SIZE && v_count < i_worm_y[7817:7812] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1303 < i_size && h_count >= i_worm_x[7823:7818] * PIXEL_SIZE && h_count < i_worm_x[7823:7818] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7823:7818] * PIXEL_SIZE && v_count < i_worm_y[7823:7818] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1304 < i_size && h_count >= i_worm_x[7829:7824] * PIXEL_SIZE && h_count < i_worm_x[7829:7824] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7829:7824] * PIXEL_SIZE && v_count < i_worm_y[7829:7824] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1305 < i_size && h_count >= i_worm_x[7835:7830] * PIXEL_SIZE && h_count < i_worm_x[7835:7830] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7835:7830] * PIXEL_SIZE && v_count < i_worm_y[7835:7830] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1306 < i_size && h_count >= i_worm_x[7841:7836] * PIXEL_SIZE && h_count < i_worm_x[7841:7836] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7841:7836] * PIXEL_SIZE && v_count < i_worm_y[7841:7836] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1307 < i_size && h_count >= i_worm_x[7847:7842] * PIXEL_SIZE && h_count < i_worm_x[7847:7842] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7847:7842] * PIXEL_SIZE && v_count < i_worm_y[7847:7842] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1308 < i_size && h_count >= i_worm_x[7853:7848] * PIXEL_SIZE && h_count < i_worm_x[7853:7848] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7853:7848] * PIXEL_SIZE && v_count < i_worm_y[7853:7848] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1309 < i_size && h_count >= i_worm_x[7859:7854] * PIXEL_SIZE && h_count < i_worm_x[7859:7854] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7859:7854] * PIXEL_SIZE && v_count < i_worm_y[7859:7854] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1310 < i_size && h_count >= i_worm_x[7865:7860] * PIXEL_SIZE && h_count < i_worm_x[7865:7860] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7865:7860] * PIXEL_SIZE && v_count < i_worm_y[7865:7860] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1311 < i_size && h_count >= i_worm_x[7871:7866] * PIXEL_SIZE && h_count < i_worm_x[7871:7866] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7871:7866] * PIXEL_SIZE && v_count < i_worm_y[7871:7866] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1312 < i_size && h_count >= i_worm_x[7877:7872] * PIXEL_SIZE && h_count < i_worm_x[7877:7872] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7877:7872] * PIXEL_SIZE && v_count < i_worm_y[7877:7872] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1313 < i_size && h_count >= i_worm_x[7883:7878] * PIXEL_SIZE && h_count < i_worm_x[7883:7878] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7883:7878] * PIXEL_SIZE && v_count < i_worm_y[7883:7878] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1314 < i_size && h_count >= i_worm_x[7889:7884] * PIXEL_SIZE && h_count < i_worm_x[7889:7884] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7889:7884] * PIXEL_SIZE && v_count < i_worm_y[7889:7884] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1315 < i_size && h_count >= i_worm_x[7895:7890] * PIXEL_SIZE && h_count < i_worm_x[7895:7890] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7895:7890] * PIXEL_SIZE && v_count < i_worm_y[7895:7890] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1316 < i_size && h_count >= i_worm_x[7901:7896] * PIXEL_SIZE && h_count < i_worm_x[7901:7896] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7901:7896] * PIXEL_SIZE && v_count < i_worm_y[7901:7896] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1317 < i_size && h_count >= i_worm_x[7907:7902] * PIXEL_SIZE && h_count < i_worm_x[7907:7902] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7907:7902] * PIXEL_SIZE && v_count < i_worm_y[7907:7902] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1318 < i_size && h_count >= i_worm_x[7913:7908] * PIXEL_SIZE && h_count < i_worm_x[7913:7908] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7913:7908] * PIXEL_SIZE && v_count < i_worm_y[7913:7908] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1319 < i_size && h_count >= i_worm_x[7919:7914] * PIXEL_SIZE && h_count < i_worm_x[7919:7914] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7919:7914] * PIXEL_SIZE && v_count < i_worm_y[7919:7914] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1320 < i_size && h_count >= i_worm_x[7925:7920] * PIXEL_SIZE && h_count < i_worm_x[7925:7920] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7925:7920] * PIXEL_SIZE && v_count < i_worm_y[7925:7920] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1321 < i_size && h_count >= i_worm_x[7931:7926] * PIXEL_SIZE && h_count < i_worm_x[7931:7926] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7931:7926] * PIXEL_SIZE && v_count < i_worm_y[7931:7926] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1322 < i_size && h_count >= i_worm_x[7937:7932] * PIXEL_SIZE && h_count < i_worm_x[7937:7932] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7937:7932] * PIXEL_SIZE && v_count < i_worm_y[7937:7932] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1323 < i_size && h_count >= i_worm_x[7943:7938] * PIXEL_SIZE && h_count < i_worm_x[7943:7938] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7943:7938] * PIXEL_SIZE && v_count < i_worm_y[7943:7938] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1324 < i_size && h_count >= i_worm_x[7949:7944] * PIXEL_SIZE && h_count < i_worm_x[7949:7944] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7949:7944] * PIXEL_SIZE && v_count < i_worm_y[7949:7944] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1325 < i_size && h_count >= i_worm_x[7955:7950] * PIXEL_SIZE && h_count < i_worm_x[7955:7950] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7955:7950] * PIXEL_SIZE && v_count < i_worm_y[7955:7950] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1326 < i_size && h_count >= i_worm_x[7961:7956] * PIXEL_SIZE && h_count < i_worm_x[7961:7956] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7961:7956] * PIXEL_SIZE && v_count < i_worm_y[7961:7956] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1327 < i_size && h_count >= i_worm_x[7967:7962] * PIXEL_SIZE && h_count < i_worm_x[7967:7962] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7967:7962] * PIXEL_SIZE && v_count < i_worm_y[7967:7962] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1328 < i_size && h_count >= i_worm_x[7973:7968] * PIXEL_SIZE && h_count < i_worm_x[7973:7968] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7973:7968] * PIXEL_SIZE && v_count < i_worm_y[7973:7968] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1329 < i_size && h_count >= i_worm_x[7979:7974] * PIXEL_SIZE && h_count < i_worm_x[7979:7974] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7979:7974] * PIXEL_SIZE && v_count < i_worm_y[7979:7974] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1330 < i_size && h_count >= i_worm_x[7985:7980] * PIXEL_SIZE && h_count < i_worm_x[7985:7980] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7985:7980] * PIXEL_SIZE && v_count < i_worm_y[7985:7980] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1331 < i_size && h_count >= i_worm_x[7991:7986] * PIXEL_SIZE && h_count < i_worm_x[7991:7986] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7991:7986] * PIXEL_SIZE && v_count < i_worm_y[7991:7986] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1332 < i_size && h_count >= i_worm_x[7997:7992] * PIXEL_SIZE && h_count < i_worm_x[7997:7992] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[7997:7992] * PIXEL_SIZE && v_count < i_worm_y[7997:7992] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1333 < i_size && h_count >= i_worm_x[8003:7998] * PIXEL_SIZE && h_count < i_worm_x[8003:7998] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8003:7998] * PIXEL_SIZE && v_count < i_worm_y[8003:7998] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1334 < i_size && h_count >= i_worm_x[8009:8004] * PIXEL_SIZE && h_count < i_worm_x[8009:8004] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8009:8004] * PIXEL_SIZE && v_count < i_worm_y[8009:8004] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1335 < i_size && h_count >= i_worm_x[8015:8010] * PIXEL_SIZE && h_count < i_worm_x[8015:8010] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8015:8010] * PIXEL_SIZE && v_count < i_worm_y[8015:8010] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1336 < i_size && h_count >= i_worm_x[8021:8016] * PIXEL_SIZE && h_count < i_worm_x[8021:8016] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8021:8016] * PIXEL_SIZE && v_count < i_worm_y[8021:8016] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1337 < i_size && h_count >= i_worm_x[8027:8022] * PIXEL_SIZE && h_count < i_worm_x[8027:8022] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8027:8022] * PIXEL_SIZE && v_count < i_worm_y[8027:8022] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1338 < i_size && h_count >= i_worm_x[8033:8028] * PIXEL_SIZE && h_count < i_worm_x[8033:8028] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8033:8028] * PIXEL_SIZE && v_count < i_worm_y[8033:8028] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1339 < i_size && h_count >= i_worm_x[8039:8034] * PIXEL_SIZE && h_count < i_worm_x[8039:8034] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8039:8034] * PIXEL_SIZE && v_count < i_worm_y[8039:8034] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1340 < i_size && h_count >= i_worm_x[8045:8040] * PIXEL_SIZE && h_count < i_worm_x[8045:8040] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8045:8040] * PIXEL_SIZE && v_count < i_worm_y[8045:8040] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1341 < i_size && h_count >= i_worm_x[8051:8046] * PIXEL_SIZE && h_count < i_worm_x[8051:8046] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8051:8046] * PIXEL_SIZE && v_count < i_worm_y[8051:8046] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1342 < i_size && h_count >= i_worm_x[8057:8052] * PIXEL_SIZE && h_count < i_worm_x[8057:8052] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8057:8052] * PIXEL_SIZE && v_count < i_worm_y[8057:8052] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1343 < i_size && h_count >= i_worm_x[8063:8058] * PIXEL_SIZE && h_count < i_worm_x[8063:8058] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8063:8058] * PIXEL_SIZE && v_count < i_worm_y[8063:8058] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1344 < i_size && h_count >= i_worm_x[8069:8064] * PIXEL_SIZE && h_count < i_worm_x[8069:8064] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8069:8064] * PIXEL_SIZE && v_count < i_worm_y[8069:8064] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1345 < i_size && h_count >= i_worm_x[8075:8070] * PIXEL_SIZE && h_count < i_worm_x[8075:8070] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8075:8070] * PIXEL_SIZE && v_count < i_worm_y[8075:8070] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1346 < i_size && h_count >= i_worm_x[8081:8076] * PIXEL_SIZE && h_count < i_worm_x[8081:8076] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8081:8076] * PIXEL_SIZE && v_count < i_worm_y[8081:8076] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1347 < i_size && h_count >= i_worm_x[8087:8082] * PIXEL_SIZE && h_count < i_worm_x[8087:8082] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8087:8082] * PIXEL_SIZE && v_count < i_worm_y[8087:8082] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1348 < i_size && h_count >= i_worm_x[8093:8088] * PIXEL_SIZE && h_count < i_worm_x[8093:8088] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8093:8088] * PIXEL_SIZE && v_count < i_worm_y[8093:8088] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1349 < i_size && h_count >= i_worm_x[8099:8094] * PIXEL_SIZE && h_count < i_worm_x[8099:8094] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8099:8094] * PIXEL_SIZE && v_count < i_worm_y[8099:8094] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1350 < i_size && h_count >= i_worm_x[8105:8100] * PIXEL_SIZE && h_count < i_worm_x[8105:8100] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8105:8100] * PIXEL_SIZE && v_count < i_worm_y[8105:8100] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1351 < i_size && h_count >= i_worm_x[8111:8106] * PIXEL_SIZE && h_count < i_worm_x[8111:8106] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8111:8106] * PIXEL_SIZE && v_count < i_worm_y[8111:8106] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1352 < i_size && h_count >= i_worm_x[8117:8112] * PIXEL_SIZE && h_count < i_worm_x[8117:8112] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8117:8112] * PIXEL_SIZE && v_count < i_worm_y[8117:8112] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1353 < i_size && h_count >= i_worm_x[8123:8118] * PIXEL_SIZE && h_count < i_worm_x[8123:8118] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8123:8118] * PIXEL_SIZE && v_count < i_worm_y[8123:8118] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1354 < i_size && h_count >= i_worm_x[8129:8124] * PIXEL_SIZE && h_count < i_worm_x[8129:8124] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8129:8124] * PIXEL_SIZE && v_count < i_worm_y[8129:8124] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1355 < i_size && h_count >= i_worm_x[8135:8130] * PIXEL_SIZE && h_count < i_worm_x[8135:8130] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8135:8130] * PIXEL_SIZE && v_count < i_worm_y[8135:8130] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1356 < i_size && h_count >= i_worm_x[8141:8136] * PIXEL_SIZE && h_count < i_worm_x[8141:8136] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8141:8136] * PIXEL_SIZE && v_count < i_worm_y[8141:8136] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1357 < i_size && h_count >= i_worm_x[8147:8142] * PIXEL_SIZE && h_count < i_worm_x[8147:8142] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8147:8142] * PIXEL_SIZE && v_count < i_worm_y[8147:8142] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1358 < i_size && h_count >= i_worm_x[8153:8148] * PIXEL_SIZE && h_count < i_worm_x[8153:8148] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8153:8148] * PIXEL_SIZE && v_count < i_worm_y[8153:8148] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1359 < i_size && h_count >= i_worm_x[8159:8154] * PIXEL_SIZE && h_count < i_worm_x[8159:8154] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8159:8154] * PIXEL_SIZE && v_count < i_worm_y[8159:8154] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1360 < i_size && h_count >= i_worm_x[8165:8160] * PIXEL_SIZE && h_count < i_worm_x[8165:8160] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8165:8160] * PIXEL_SIZE && v_count < i_worm_y[8165:8160] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1361 < i_size && h_count >= i_worm_x[8171:8166] * PIXEL_SIZE && h_count < i_worm_x[8171:8166] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8171:8166] * PIXEL_SIZE && v_count < i_worm_y[8171:8166] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1362 < i_size && h_count >= i_worm_x[8177:8172] * PIXEL_SIZE && h_count < i_worm_x[8177:8172] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8177:8172] * PIXEL_SIZE && v_count < i_worm_y[8177:8172] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1363 < i_size && h_count >= i_worm_x[8183:8178] * PIXEL_SIZE && h_count < i_worm_x[8183:8178] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8183:8178] * PIXEL_SIZE && v_count < i_worm_y[8183:8178] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1364 < i_size && h_count >= i_worm_x[8189:8184] * PIXEL_SIZE && h_count < i_worm_x[8189:8184] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8189:8184] * PIXEL_SIZE && v_count < i_worm_y[8189:8184] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1365 < i_size && h_count >= i_worm_x[8195:8190] * PIXEL_SIZE && h_count < i_worm_x[8195:8190] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8195:8190] * PIXEL_SIZE && v_count < i_worm_y[8195:8190] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1366 < i_size && h_count >= i_worm_x[8201:8196] * PIXEL_SIZE && h_count < i_worm_x[8201:8196] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8201:8196] * PIXEL_SIZE && v_count < i_worm_y[8201:8196] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1367 < i_size && h_count >= i_worm_x[8207:8202] * PIXEL_SIZE && h_count < i_worm_x[8207:8202] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8207:8202] * PIXEL_SIZE && v_count < i_worm_y[8207:8202] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1368 < i_size && h_count >= i_worm_x[8213:8208] * PIXEL_SIZE && h_count < i_worm_x[8213:8208] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8213:8208] * PIXEL_SIZE && v_count < i_worm_y[8213:8208] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1369 < i_size && h_count >= i_worm_x[8219:8214] * PIXEL_SIZE && h_count < i_worm_x[8219:8214] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8219:8214] * PIXEL_SIZE && v_count < i_worm_y[8219:8214] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1370 < i_size && h_count >= i_worm_x[8225:8220] * PIXEL_SIZE && h_count < i_worm_x[8225:8220] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8225:8220] * PIXEL_SIZE && v_count < i_worm_y[8225:8220] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1371 < i_size && h_count >= i_worm_x[8231:8226] * PIXEL_SIZE && h_count < i_worm_x[8231:8226] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8231:8226] * PIXEL_SIZE && v_count < i_worm_y[8231:8226] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1372 < i_size && h_count >= i_worm_x[8237:8232] * PIXEL_SIZE && h_count < i_worm_x[8237:8232] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8237:8232] * PIXEL_SIZE && v_count < i_worm_y[8237:8232] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1373 < i_size && h_count >= i_worm_x[8243:8238] * PIXEL_SIZE && h_count < i_worm_x[8243:8238] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8243:8238] * PIXEL_SIZE && v_count < i_worm_y[8243:8238] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1374 < i_size && h_count >= i_worm_x[8249:8244] * PIXEL_SIZE && h_count < i_worm_x[8249:8244] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8249:8244] * PIXEL_SIZE && v_count < i_worm_y[8249:8244] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1375 < i_size && h_count >= i_worm_x[8255:8250] * PIXEL_SIZE && h_count < i_worm_x[8255:8250] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8255:8250] * PIXEL_SIZE && v_count < i_worm_y[8255:8250] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1376 < i_size && h_count >= i_worm_x[8261:8256] * PIXEL_SIZE && h_count < i_worm_x[8261:8256] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8261:8256] * PIXEL_SIZE && v_count < i_worm_y[8261:8256] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1377 < i_size && h_count >= i_worm_x[8267:8262] * PIXEL_SIZE && h_count < i_worm_x[8267:8262] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8267:8262] * PIXEL_SIZE && v_count < i_worm_y[8267:8262] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1378 < i_size && h_count >= i_worm_x[8273:8268] * PIXEL_SIZE && h_count < i_worm_x[8273:8268] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8273:8268] * PIXEL_SIZE && v_count < i_worm_y[8273:8268] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1379 < i_size && h_count >= i_worm_x[8279:8274] * PIXEL_SIZE && h_count < i_worm_x[8279:8274] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8279:8274] * PIXEL_SIZE && v_count < i_worm_y[8279:8274] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1380 < i_size && h_count >= i_worm_x[8285:8280] * PIXEL_SIZE && h_count < i_worm_x[8285:8280] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8285:8280] * PIXEL_SIZE && v_count < i_worm_y[8285:8280] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1381 < i_size && h_count >= i_worm_x[8291:8286] * PIXEL_SIZE && h_count < i_worm_x[8291:8286] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8291:8286] * PIXEL_SIZE && v_count < i_worm_y[8291:8286] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1382 < i_size && h_count >= i_worm_x[8297:8292] * PIXEL_SIZE && h_count < i_worm_x[8297:8292] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8297:8292] * PIXEL_SIZE && v_count < i_worm_y[8297:8292] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1383 < i_size && h_count >= i_worm_x[8303:8298] * PIXEL_SIZE && h_count < i_worm_x[8303:8298] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8303:8298] * PIXEL_SIZE && v_count < i_worm_y[8303:8298] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1384 < i_size && h_count >= i_worm_x[8309:8304] * PIXEL_SIZE && h_count < i_worm_x[8309:8304] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8309:8304] * PIXEL_SIZE && v_count < i_worm_y[8309:8304] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1385 < i_size && h_count >= i_worm_x[8315:8310] * PIXEL_SIZE && h_count < i_worm_x[8315:8310] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8315:8310] * PIXEL_SIZE && v_count < i_worm_y[8315:8310] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1386 < i_size && h_count >= i_worm_x[8321:8316] * PIXEL_SIZE && h_count < i_worm_x[8321:8316] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8321:8316] * PIXEL_SIZE && v_count < i_worm_y[8321:8316] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1387 < i_size && h_count >= i_worm_x[8327:8322] * PIXEL_SIZE && h_count < i_worm_x[8327:8322] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8327:8322] * PIXEL_SIZE && v_count < i_worm_y[8327:8322] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1388 < i_size && h_count >= i_worm_x[8333:8328] * PIXEL_SIZE && h_count < i_worm_x[8333:8328] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8333:8328] * PIXEL_SIZE && v_count < i_worm_y[8333:8328] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1389 < i_size && h_count >= i_worm_x[8339:8334] * PIXEL_SIZE && h_count < i_worm_x[8339:8334] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8339:8334] * PIXEL_SIZE && v_count < i_worm_y[8339:8334] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1390 < i_size && h_count >= i_worm_x[8345:8340] * PIXEL_SIZE && h_count < i_worm_x[8345:8340] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8345:8340] * PIXEL_SIZE && v_count < i_worm_y[8345:8340] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1391 < i_size && h_count >= i_worm_x[8351:8346] * PIXEL_SIZE && h_count < i_worm_x[8351:8346] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8351:8346] * PIXEL_SIZE && v_count < i_worm_y[8351:8346] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1392 < i_size && h_count >= i_worm_x[8357:8352] * PIXEL_SIZE && h_count < i_worm_x[8357:8352] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8357:8352] * PIXEL_SIZE && v_count < i_worm_y[8357:8352] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1393 < i_size && h_count >= i_worm_x[8363:8358] * PIXEL_SIZE && h_count < i_worm_x[8363:8358] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8363:8358] * PIXEL_SIZE && v_count < i_worm_y[8363:8358] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1394 < i_size && h_count >= i_worm_x[8369:8364] * PIXEL_SIZE && h_count < i_worm_x[8369:8364] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8369:8364] * PIXEL_SIZE && v_count < i_worm_y[8369:8364] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1395 < i_size && h_count >= i_worm_x[8375:8370] * PIXEL_SIZE && h_count < i_worm_x[8375:8370] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8375:8370] * PIXEL_SIZE && v_count < i_worm_y[8375:8370] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1396 < i_size && h_count >= i_worm_x[8381:8376] * PIXEL_SIZE && h_count < i_worm_x[8381:8376] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8381:8376] * PIXEL_SIZE && v_count < i_worm_y[8381:8376] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1397 < i_size && h_count >= i_worm_x[8387:8382] * PIXEL_SIZE && h_count < i_worm_x[8387:8382] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8387:8382] * PIXEL_SIZE && v_count < i_worm_y[8387:8382] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1398 < i_size && h_count >= i_worm_x[8393:8388] * PIXEL_SIZE && h_count < i_worm_x[8393:8388] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8393:8388] * PIXEL_SIZE && v_count < i_worm_y[8393:8388] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1399 < i_size && h_count >= i_worm_x[8399:8394] * PIXEL_SIZE && h_count < i_worm_x[8399:8394] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8399:8394] * PIXEL_SIZE && v_count < i_worm_y[8399:8394] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1400 < i_size && h_count >= i_worm_x[8405:8400] * PIXEL_SIZE && h_count < i_worm_x[8405:8400] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8405:8400] * PIXEL_SIZE && v_count < i_worm_y[8405:8400] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1401 < i_size && h_count >= i_worm_x[8411:8406] * PIXEL_SIZE && h_count < i_worm_x[8411:8406] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8411:8406] * PIXEL_SIZE && v_count < i_worm_y[8411:8406] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1402 < i_size && h_count >= i_worm_x[8417:8412] * PIXEL_SIZE && h_count < i_worm_x[8417:8412] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8417:8412] * PIXEL_SIZE && v_count < i_worm_y[8417:8412] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1403 < i_size && h_count >= i_worm_x[8423:8418] * PIXEL_SIZE && h_count < i_worm_x[8423:8418] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8423:8418] * PIXEL_SIZE && v_count < i_worm_y[8423:8418] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1404 < i_size && h_count >= i_worm_x[8429:8424] * PIXEL_SIZE && h_count < i_worm_x[8429:8424] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8429:8424] * PIXEL_SIZE && v_count < i_worm_y[8429:8424] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1405 < i_size && h_count >= i_worm_x[8435:8430] * PIXEL_SIZE && h_count < i_worm_x[8435:8430] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8435:8430] * PIXEL_SIZE && v_count < i_worm_y[8435:8430] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1406 < i_size && h_count >= i_worm_x[8441:8436] * PIXEL_SIZE && h_count < i_worm_x[8441:8436] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8441:8436] * PIXEL_SIZE && v_count < i_worm_y[8441:8436] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1407 < i_size && h_count >= i_worm_x[8447:8442] * PIXEL_SIZE && h_count < i_worm_x[8447:8442] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8447:8442] * PIXEL_SIZE && v_count < i_worm_y[8447:8442] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1408 < i_size && h_count >= i_worm_x[8453:8448] * PIXEL_SIZE && h_count < i_worm_x[8453:8448] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8453:8448] * PIXEL_SIZE && v_count < i_worm_y[8453:8448] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1409 < i_size && h_count >= i_worm_x[8459:8454] * PIXEL_SIZE && h_count < i_worm_x[8459:8454] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8459:8454] * PIXEL_SIZE && v_count < i_worm_y[8459:8454] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1410 < i_size && h_count >= i_worm_x[8465:8460] * PIXEL_SIZE && h_count < i_worm_x[8465:8460] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8465:8460] * PIXEL_SIZE && v_count < i_worm_y[8465:8460] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1411 < i_size && h_count >= i_worm_x[8471:8466] * PIXEL_SIZE && h_count < i_worm_x[8471:8466] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8471:8466] * PIXEL_SIZE && v_count < i_worm_y[8471:8466] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1412 < i_size && h_count >= i_worm_x[8477:8472] * PIXEL_SIZE && h_count < i_worm_x[8477:8472] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8477:8472] * PIXEL_SIZE && v_count < i_worm_y[8477:8472] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1413 < i_size && h_count >= i_worm_x[8483:8478] * PIXEL_SIZE && h_count < i_worm_x[8483:8478] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8483:8478] * PIXEL_SIZE && v_count < i_worm_y[8483:8478] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1414 < i_size && h_count >= i_worm_x[8489:8484] * PIXEL_SIZE && h_count < i_worm_x[8489:8484] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8489:8484] * PIXEL_SIZE && v_count < i_worm_y[8489:8484] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1415 < i_size && h_count >= i_worm_x[8495:8490] * PIXEL_SIZE && h_count < i_worm_x[8495:8490] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8495:8490] * PIXEL_SIZE && v_count < i_worm_y[8495:8490] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1416 < i_size && h_count >= i_worm_x[8501:8496] * PIXEL_SIZE && h_count < i_worm_x[8501:8496] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8501:8496] * PIXEL_SIZE && v_count < i_worm_y[8501:8496] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1417 < i_size && h_count >= i_worm_x[8507:8502] * PIXEL_SIZE && h_count < i_worm_x[8507:8502] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8507:8502] * PIXEL_SIZE && v_count < i_worm_y[8507:8502] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1418 < i_size && h_count >= i_worm_x[8513:8508] * PIXEL_SIZE && h_count < i_worm_x[8513:8508] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8513:8508] * PIXEL_SIZE && v_count < i_worm_y[8513:8508] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1419 < i_size && h_count >= i_worm_x[8519:8514] * PIXEL_SIZE && h_count < i_worm_x[8519:8514] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8519:8514] * PIXEL_SIZE && v_count < i_worm_y[8519:8514] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1420 < i_size && h_count >= i_worm_x[8525:8520] * PIXEL_SIZE && h_count < i_worm_x[8525:8520] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8525:8520] * PIXEL_SIZE && v_count < i_worm_y[8525:8520] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1421 < i_size && h_count >= i_worm_x[8531:8526] * PIXEL_SIZE && h_count < i_worm_x[8531:8526] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8531:8526] * PIXEL_SIZE && v_count < i_worm_y[8531:8526] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1422 < i_size && h_count >= i_worm_x[8537:8532] * PIXEL_SIZE && h_count < i_worm_x[8537:8532] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8537:8532] * PIXEL_SIZE && v_count < i_worm_y[8537:8532] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1423 < i_size && h_count >= i_worm_x[8543:8538] * PIXEL_SIZE && h_count < i_worm_x[8543:8538] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8543:8538] * PIXEL_SIZE && v_count < i_worm_y[8543:8538] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1424 < i_size && h_count >= i_worm_x[8549:8544] * PIXEL_SIZE && h_count < i_worm_x[8549:8544] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8549:8544] * PIXEL_SIZE && v_count < i_worm_y[8549:8544] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1425 < i_size && h_count >= i_worm_x[8555:8550] * PIXEL_SIZE && h_count < i_worm_x[8555:8550] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8555:8550] * PIXEL_SIZE && v_count < i_worm_y[8555:8550] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1426 < i_size && h_count >= i_worm_x[8561:8556] * PIXEL_SIZE && h_count < i_worm_x[8561:8556] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8561:8556] * PIXEL_SIZE && v_count < i_worm_y[8561:8556] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1427 < i_size && h_count >= i_worm_x[8567:8562] * PIXEL_SIZE && h_count < i_worm_x[8567:8562] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8567:8562] * PIXEL_SIZE && v_count < i_worm_y[8567:8562] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1428 < i_size && h_count >= i_worm_x[8573:8568] * PIXEL_SIZE && h_count < i_worm_x[8573:8568] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8573:8568] * PIXEL_SIZE && v_count < i_worm_y[8573:8568] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1429 < i_size && h_count >= i_worm_x[8579:8574] * PIXEL_SIZE && h_count < i_worm_x[8579:8574] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8579:8574] * PIXEL_SIZE && v_count < i_worm_y[8579:8574] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1430 < i_size && h_count >= i_worm_x[8585:8580] * PIXEL_SIZE && h_count < i_worm_x[8585:8580] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8585:8580] * PIXEL_SIZE && v_count < i_worm_y[8585:8580] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1431 < i_size && h_count >= i_worm_x[8591:8586] * PIXEL_SIZE && h_count < i_worm_x[8591:8586] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8591:8586] * PIXEL_SIZE && v_count < i_worm_y[8591:8586] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1432 < i_size && h_count >= i_worm_x[8597:8592] * PIXEL_SIZE && h_count < i_worm_x[8597:8592] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8597:8592] * PIXEL_SIZE && v_count < i_worm_y[8597:8592] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1433 < i_size && h_count >= i_worm_x[8603:8598] * PIXEL_SIZE && h_count < i_worm_x[8603:8598] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8603:8598] * PIXEL_SIZE && v_count < i_worm_y[8603:8598] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1434 < i_size && h_count >= i_worm_x[8609:8604] * PIXEL_SIZE && h_count < i_worm_x[8609:8604] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8609:8604] * PIXEL_SIZE && v_count < i_worm_y[8609:8604] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1435 < i_size && h_count >= i_worm_x[8615:8610] * PIXEL_SIZE && h_count < i_worm_x[8615:8610] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8615:8610] * PIXEL_SIZE && v_count < i_worm_y[8615:8610] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1436 < i_size && h_count >= i_worm_x[8621:8616] * PIXEL_SIZE && h_count < i_worm_x[8621:8616] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8621:8616] * PIXEL_SIZE && v_count < i_worm_y[8621:8616] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1437 < i_size && h_count >= i_worm_x[8627:8622] * PIXEL_SIZE && h_count < i_worm_x[8627:8622] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8627:8622] * PIXEL_SIZE && v_count < i_worm_y[8627:8622] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1438 < i_size && h_count >= i_worm_x[8633:8628] * PIXEL_SIZE && h_count < i_worm_x[8633:8628] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8633:8628] * PIXEL_SIZE && v_count < i_worm_y[8633:8628] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1439 < i_size && h_count >= i_worm_x[8639:8634] * PIXEL_SIZE && h_count < i_worm_x[8639:8634] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8639:8634] * PIXEL_SIZE && v_count < i_worm_y[8639:8634] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1440 < i_size && h_count >= i_worm_x[8645:8640] * PIXEL_SIZE && h_count < i_worm_x[8645:8640] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8645:8640] * PIXEL_SIZE && v_count < i_worm_y[8645:8640] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1441 < i_size && h_count >= i_worm_x[8651:8646] * PIXEL_SIZE && h_count < i_worm_x[8651:8646] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8651:8646] * PIXEL_SIZE && v_count < i_worm_y[8651:8646] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1442 < i_size && h_count >= i_worm_x[8657:8652] * PIXEL_SIZE && h_count < i_worm_x[8657:8652] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8657:8652] * PIXEL_SIZE && v_count < i_worm_y[8657:8652] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1443 < i_size && h_count >= i_worm_x[8663:8658] * PIXEL_SIZE && h_count < i_worm_x[8663:8658] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8663:8658] * PIXEL_SIZE && v_count < i_worm_y[8663:8658] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1444 < i_size && h_count >= i_worm_x[8669:8664] * PIXEL_SIZE && h_count < i_worm_x[8669:8664] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8669:8664] * PIXEL_SIZE && v_count < i_worm_y[8669:8664] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1445 < i_size && h_count >= i_worm_x[8675:8670] * PIXEL_SIZE && h_count < i_worm_x[8675:8670] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8675:8670] * PIXEL_SIZE && v_count < i_worm_y[8675:8670] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1446 < i_size && h_count >= i_worm_x[8681:8676] * PIXEL_SIZE && h_count < i_worm_x[8681:8676] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8681:8676] * PIXEL_SIZE && v_count < i_worm_y[8681:8676] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1447 < i_size && h_count >= i_worm_x[8687:8682] * PIXEL_SIZE && h_count < i_worm_x[8687:8682] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8687:8682] * PIXEL_SIZE && v_count < i_worm_y[8687:8682] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1448 < i_size && h_count >= i_worm_x[8693:8688] * PIXEL_SIZE && h_count < i_worm_x[8693:8688] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8693:8688] * PIXEL_SIZE && v_count < i_worm_y[8693:8688] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1449 < i_size && h_count >= i_worm_x[8699:8694] * PIXEL_SIZE && h_count < i_worm_x[8699:8694] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8699:8694] * PIXEL_SIZE && v_count < i_worm_y[8699:8694] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1450 < i_size && h_count >= i_worm_x[8705:8700] * PIXEL_SIZE && h_count < i_worm_x[8705:8700] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8705:8700] * PIXEL_SIZE && v_count < i_worm_y[8705:8700] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1451 < i_size && h_count >= i_worm_x[8711:8706] * PIXEL_SIZE && h_count < i_worm_x[8711:8706] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8711:8706] * PIXEL_SIZE && v_count < i_worm_y[8711:8706] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1452 < i_size && h_count >= i_worm_x[8717:8712] * PIXEL_SIZE && h_count < i_worm_x[8717:8712] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8717:8712] * PIXEL_SIZE && v_count < i_worm_y[8717:8712] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1453 < i_size && h_count >= i_worm_x[8723:8718] * PIXEL_SIZE && h_count < i_worm_x[8723:8718] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8723:8718] * PIXEL_SIZE && v_count < i_worm_y[8723:8718] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1454 < i_size && h_count >= i_worm_x[8729:8724] * PIXEL_SIZE && h_count < i_worm_x[8729:8724] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8729:8724] * PIXEL_SIZE && v_count < i_worm_y[8729:8724] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1455 < i_size && h_count >= i_worm_x[8735:8730] * PIXEL_SIZE && h_count < i_worm_x[8735:8730] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8735:8730] * PIXEL_SIZE && v_count < i_worm_y[8735:8730] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1456 < i_size && h_count >= i_worm_x[8741:8736] * PIXEL_SIZE && h_count < i_worm_x[8741:8736] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8741:8736] * PIXEL_SIZE && v_count < i_worm_y[8741:8736] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1457 < i_size && h_count >= i_worm_x[8747:8742] * PIXEL_SIZE && h_count < i_worm_x[8747:8742] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8747:8742] * PIXEL_SIZE && v_count < i_worm_y[8747:8742] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1458 < i_size && h_count >= i_worm_x[8753:8748] * PIXEL_SIZE && h_count < i_worm_x[8753:8748] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8753:8748] * PIXEL_SIZE && v_count < i_worm_y[8753:8748] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1459 < i_size && h_count >= i_worm_x[8759:8754] * PIXEL_SIZE && h_count < i_worm_x[8759:8754] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8759:8754] * PIXEL_SIZE && v_count < i_worm_y[8759:8754] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1460 < i_size && h_count >= i_worm_x[8765:8760] * PIXEL_SIZE && h_count < i_worm_x[8765:8760] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8765:8760] * PIXEL_SIZE && v_count < i_worm_y[8765:8760] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1461 < i_size && h_count >= i_worm_x[8771:8766] * PIXEL_SIZE && h_count < i_worm_x[8771:8766] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8771:8766] * PIXEL_SIZE && v_count < i_worm_y[8771:8766] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1462 < i_size && h_count >= i_worm_x[8777:8772] * PIXEL_SIZE && h_count < i_worm_x[8777:8772] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8777:8772] * PIXEL_SIZE && v_count < i_worm_y[8777:8772] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1463 < i_size && h_count >= i_worm_x[8783:8778] * PIXEL_SIZE && h_count < i_worm_x[8783:8778] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8783:8778] * PIXEL_SIZE && v_count < i_worm_y[8783:8778] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1464 < i_size && h_count >= i_worm_x[8789:8784] * PIXEL_SIZE && h_count < i_worm_x[8789:8784] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8789:8784] * PIXEL_SIZE && v_count < i_worm_y[8789:8784] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1465 < i_size && h_count >= i_worm_x[8795:8790] * PIXEL_SIZE && h_count < i_worm_x[8795:8790] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8795:8790] * PIXEL_SIZE && v_count < i_worm_y[8795:8790] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1466 < i_size && h_count >= i_worm_x[8801:8796] * PIXEL_SIZE && h_count < i_worm_x[8801:8796] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8801:8796] * PIXEL_SIZE && v_count < i_worm_y[8801:8796] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1467 < i_size && h_count >= i_worm_x[8807:8802] * PIXEL_SIZE && h_count < i_worm_x[8807:8802] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8807:8802] * PIXEL_SIZE && v_count < i_worm_y[8807:8802] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1468 < i_size && h_count >= i_worm_x[8813:8808] * PIXEL_SIZE && h_count < i_worm_x[8813:8808] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8813:8808] * PIXEL_SIZE && v_count < i_worm_y[8813:8808] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1469 < i_size && h_count >= i_worm_x[8819:8814] * PIXEL_SIZE && h_count < i_worm_x[8819:8814] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8819:8814] * PIXEL_SIZE && v_count < i_worm_y[8819:8814] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1470 < i_size && h_count >= i_worm_x[8825:8820] * PIXEL_SIZE && h_count < i_worm_x[8825:8820] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8825:8820] * PIXEL_SIZE && v_count < i_worm_y[8825:8820] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1471 < i_size && h_count >= i_worm_x[8831:8826] * PIXEL_SIZE && h_count < i_worm_x[8831:8826] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8831:8826] * PIXEL_SIZE && v_count < i_worm_y[8831:8826] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1472 < i_size && h_count >= i_worm_x[8837:8832] * PIXEL_SIZE && h_count < i_worm_x[8837:8832] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8837:8832] * PIXEL_SIZE && v_count < i_worm_y[8837:8832] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1473 < i_size && h_count >= i_worm_x[8843:8838] * PIXEL_SIZE && h_count < i_worm_x[8843:8838] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8843:8838] * PIXEL_SIZE && v_count < i_worm_y[8843:8838] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1474 < i_size && h_count >= i_worm_x[8849:8844] * PIXEL_SIZE && h_count < i_worm_x[8849:8844] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8849:8844] * PIXEL_SIZE && v_count < i_worm_y[8849:8844] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1475 < i_size && h_count >= i_worm_x[8855:8850] * PIXEL_SIZE && h_count < i_worm_x[8855:8850] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8855:8850] * PIXEL_SIZE && v_count < i_worm_y[8855:8850] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1476 < i_size && h_count >= i_worm_x[8861:8856] * PIXEL_SIZE && h_count < i_worm_x[8861:8856] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8861:8856] * PIXEL_SIZE && v_count < i_worm_y[8861:8856] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1477 < i_size && h_count >= i_worm_x[8867:8862] * PIXEL_SIZE && h_count < i_worm_x[8867:8862] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8867:8862] * PIXEL_SIZE && v_count < i_worm_y[8867:8862] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1478 < i_size && h_count >= i_worm_x[8873:8868] * PIXEL_SIZE && h_count < i_worm_x[8873:8868] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8873:8868] * PIXEL_SIZE && v_count < i_worm_y[8873:8868] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1479 < i_size && h_count >= i_worm_x[8879:8874] * PIXEL_SIZE && h_count < i_worm_x[8879:8874] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8879:8874] * PIXEL_SIZE && v_count < i_worm_y[8879:8874] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1480 < i_size && h_count >= i_worm_x[8885:8880] * PIXEL_SIZE && h_count < i_worm_x[8885:8880] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8885:8880] * PIXEL_SIZE && v_count < i_worm_y[8885:8880] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1481 < i_size && h_count >= i_worm_x[8891:8886] * PIXEL_SIZE && h_count < i_worm_x[8891:8886] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8891:8886] * PIXEL_SIZE && v_count < i_worm_y[8891:8886] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1482 < i_size && h_count >= i_worm_x[8897:8892] * PIXEL_SIZE && h_count < i_worm_x[8897:8892] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8897:8892] * PIXEL_SIZE && v_count < i_worm_y[8897:8892] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1483 < i_size && h_count >= i_worm_x[8903:8898] * PIXEL_SIZE && h_count < i_worm_x[8903:8898] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8903:8898] * PIXEL_SIZE && v_count < i_worm_y[8903:8898] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1484 < i_size && h_count >= i_worm_x[8909:8904] * PIXEL_SIZE && h_count < i_worm_x[8909:8904] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8909:8904] * PIXEL_SIZE && v_count < i_worm_y[8909:8904] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1485 < i_size && h_count >= i_worm_x[8915:8910] * PIXEL_SIZE && h_count < i_worm_x[8915:8910] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8915:8910] * PIXEL_SIZE && v_count < i_worm_y[8915:8910] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1486 < i_size && h_count >= i_worm_x[8921:8916] * PIXEL_SIZE && h_count < i_worm_x[8921:8916] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8921:8916] * PIXEL_SIZE && v_count < i_worm_y[8921:8916] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1487 < i_size && h_count >= i_worm_x[8927:8922] * PIXEL_SIZE && h_count < i_worm_x[8927:8922] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8927:8922] * PIXEL_SIZE && v_count < i_worm_y[8927:8922] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1488 < i_size && h_count >= i_worm_x[8933:8928] * PIXEL_SIZE && h_count < i_worm_x[8933:8928] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8933:8928] * PIXEL_SIZE && v_count < i_worm_y[8933:8928] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1489 < i_size && h_count >= i_worm_x[8939:8934] * PIXEL_SIZE && h_count < i_worm_x[8939:8934] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8939:8934] * PIXEL_SIZE && v_count < i_worm_y[8939:8934] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1490 < i_size && h_count >= i_worm_x[8945:8940] * PIXEL_SIZE && h_count < i_worm_x[8945:8940] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8945:8940] * PIXEL_SIZE && v_count < i_worm_y[8945:8940] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1491 < i_size && h_count >= i_worm_x[8951:8946] * PIXEL_SIZE && h_count < i_worm_x[8951:8946] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8951:8946] * PIXEL_SIZE && v_count < i_worm_y[8951:8946] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1492 < i_size && h_count >= i_worm_x[8957:8952] * PIXEL_SIZE && h_count < i_worm_x[8957:8952] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8957:8952] * PIXEL_SIZE && v_count < i_worm_y[8957:8952] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1493 < i_size && h_count >= i_worm_x[8963:8958] * PIXEL_SIZE && h_count < i_worm_x[8963:8958] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8963:8958] * PIXEL_SIZE && v_count < i_worm_y[8963:8958] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1494 < i_size && h_count >= i_worm_x[8969:8964] * PIXEL_SIZE && h_count < i_worm_x[8969:8964] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8969:8964] * PIXEL_SIZE && v_count < i_worm_y[8969:8964] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1495 < i_size && h_count >= i_worm_x[8975:8970] * PIXEL_SIZE && h_count < i_worm_x[8975:8970] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8975:8970] * PIXEL_SIZE && v_count < i_worm_y[8975:8970] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1496 < i_size && h_count >= i_worm_x[8981:8976] * PIXEL_SIZE && h_count < i_worm_x[8981:8976] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8981:8976] * PIXEL_SIZE && v_count < i_worm_y[8981:8976] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1497 < i_size && h_count >= i_worm_x[8987:8982] * PIXEL_SIZE && h_count < i_worm_x[8987:8982] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8987:8982] * PIXEL_SIZE && v_count < i_worm_y[8987:8982] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1498 < i_size && h_count >= i_worm_x[8993:8988] * PIXEL_SIZE && h_count < i_worm_x[8993:8988] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8993:8988] * PIXEL_SIZE && v_count < i_worm_y[8993:8988] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1499 < i_size && h_count >= i_worm_x[8999:8994] * PIXEL_SIZE && h_count < i_worm_x[8999:8994] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[8999:8994] * PIXEL_SIZE && v_count < i_worm_y[8999:8994] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1500 < i_size && h_count >= i_worm_x[9005:9000] * PIXEL_SIZE && h_count < i_worm_x[9005:9000] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9005:9000] * PIXEL_SIZE && v_count < i_worm_y[9005:9000] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1501 < i_size && h_count >= i_worm_x[9011:9006] * PIXEL_SIZE && h_count < i_worm_x[9011:9006] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9011:9006] * PIXEL_SIZE && v_count < i_worm_y[9011:9006] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1502 < i_size && h_count >= i_worm_x[9017:9012] * PIXEL_SIZE && h_count < i_worm_x[9017:9012] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9017:9012] * PIXEL_SIZE && v_count < i_worm_y[9017:9012] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1503 < i_size && h_count >= i_worm_x[9023:9018] * PIXEL_SIZE && h_count < i_worm_x[9023:9018] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9023:9018] * PIXEL_SIZE && v_count < i_worm_y[9023:9018] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1504 < i_size && h_count >= i_worm_x[9029:9024] * PIXEL_SIZE && h_count < i_worm_x[9029:9024] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9029:9024] * PIXEL_SIZE && v_count < i_worm_y[9029:9024] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1505 < i_size && h_count >= i_worm_x[9035:9030] * PIXEL_SIZE && h_count < i_worm_x[9035:9030] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9035:9030] * PIXEL_SIZE && v_count < i_worm_y[9035:9030] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1506 < i_size && h_count >= i_worm_x[9041:9036] * PIXEL_SIZE && h_count < i_worm_x[9041:9036] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9041:9036] * PIXEL_SIZE && v_count < i_worm_y[9041:9036] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1507 < i_size && h_count >= i_worm_x[9047:9042] * PIXEL_SIZE && h_count < i_worm_x[9047:9042] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9047:9042] * PIXEL_SIZE && v_count < i_worm_y[9047:9042] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1508 < i_size && h_count >= i_worm_x[9053:9048] * PIXEL_SIZE && h_count < i_worm_x[9053:9048] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9053:9048] * PIXEL_SIZE && v_count < i_worm_y[9053:9048] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1509 < i_size && h_count >= i_worm_x[9059:9054] * PIXEL_SIZE && h_count < i_worm_x[9059:9054] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9059:9054] * PIXEL_SIZE && v_count < i_worm_y[9059:9054] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1510 < i_size && h_count >= i_worm_x[9065:9060] * PIXEL_SIZE && h_count < i_worm_x[9065:9060] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9065:9060] * PIXEL_SIZE && v_count < i_worm_y[9065:9060] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1511 < i_size && h_count >= i_worm_x[9071:9066] * PIXEL_SIZE && h_count < i_worm_x[9071:9066] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9071:9066] * PIXEL_SIZE && v_count < i_worm_y[9071:9066] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1512 < i_size && h_count >= i_worm_x[9077:9072] * PIXEL_SIZE && h_count < i_worm_x[9077:9072] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9077:9072] * PIXEL_SIZE && v_count < i_worm_y[9077:9072] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1513 < i_size && h_count >= i_worm_x[9083:9078] * PIXEL_SIZE && h_count < i_worm_x[9083:9078] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9083:9078] * PIXEL_SIZE && v_count < i_worm_y[9083:9078] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1514 < i_size && h_count >= i_worm_x[9089:9084] * PIXEL_SIZE && h_count < i_worm_x[9089:9084] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9089:9084] * PIXEL_SIZE && v_count < i_worm_y[9089:9084] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1515 < i_size && h_count >= i_worm_x[9095:9090] * PIXEL_SIZE && h_count < i_worm_x[9095:9090] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9095:9090] * PIXEL_SIZE && v_count < i_worm_y[9095:9090] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1516 < i_size && h_count >= i_worm_x[9101:9096] * PIXEL_SIZE && h_count < i_worm_x[9101:9096] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9101:9096] * PIXEL_SIZE && v_count < i_worm_y[9101:9096] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1517 < i_size && h_count >= i_worm_x[9107:9102] * PIXEL_SIZE && h_count < i_worm_x[9107:9102] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9107:9102] * PIXEL_SIZE && v_count < i_worm_y[9107:9102] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1518 < i_size && h_count >= i_worm_x[9113:9108] * PIXEL_SIZE && h_count < i_worm_x[9113:9108] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9113:9108] * PIXEL_SIZE && v_count < i_worm_y[9113:9108] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1519 < i_size && h_count >= i_worm_x[9119:9114] * PIXEL_SIZE && h_count < i_worm_x[9119:9114] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9119:9114] * PIXEL_SIZE && v_count < i_worm_y[9119:9114] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1520 < i_size && h_count >= i_worm_x[9125:9120] * PIXEL_SIZE && h_count < i_worm_x[9125:9120] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9125:9120] * PIXEL_SIZE && v_count < i_worm_y[9125:9120] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1521 < i_size && h_count >= i_worm_x[9131:9126] * PIXEL_SIZE && h_count < i_worm_x[9131:9126] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9131:9126] * PIXEL_SIZE && v_count < i_worm_y[9131:9126] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1522 < i_size && h_count >= i_worm_x[9137:9132] * PIXEL_SIZE && h_count < i_worm_x[9137:9132] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9137:9132] * PIXEL_SIZE && v_count < i_worm_y[9137:9132] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1523 < i_size && h_count >= i_worm_x[9143:9138] * PIXEL_SIZE && h_count < i_worm_x[9143:9138] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9143:9138] * PIXEL_SIZE && v_count < i_worm_y[9143:9138] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1524 < i_size && h_count >= i_worm_x[9149:9144] * PIXEL_SIZE && h_count < i_worm_x[9149:9144] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9149:9144] * PIXEL_SIZE && v_count < i_worm_y[9149:9144] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1525 < i_size && h_count >= i_worm_x[9155:9150] * PIXEL_SIZE && h_count < i_worm_x[9155:9150] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9155:9150] * PIXEL_SIZE && v_count < i_worm_y[9155:9150] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1526 < i_size && h_count >= i_worm_x[9161:9156] * PIXEL_SIZE && h_count < i_worm_x[9161:9156] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9161:9156] * PIXEL_SIZE && v_count < i_worm_y[9161:9156] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1527 < i_size && h_count >= i_worm_x[9167:9162] * PIXEL_SIZE && h_count < i_worm_x[9167:9162] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9167:9162] * PIXEL_SIZE && v_count < i_worm_y[9167:9162] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1528 < i_size && h_count >= i_worm_x[9173:9168] * PIXEL_SIZE && h_count < i_worm_x[9173:9168] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9173:9168] * PIXEL_SIZE && v_count < i_worm_y[9173:9168] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1529 < i_size && h_count >= i_worm_x[9179:9174] * PIXEL_SIZE && h_count < i_worm_x[9179:9174] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9179:9174] * PIXEL_SIZE && v_count < i_worm_y[9179:9174] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1530 < i_size && h_count >= i_worm_x[9185:9180] * PIXEL_SIZE && h_count < i_worm_x[9185:9180] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9185:9180] * PIXEL_SIZE && v_count < i_worm_y[9185:9180] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1531 < i_size && h_count >= i_worm_x[9191:9186] * PIXEL_SIZE && h_count < i_worm_x[9191:9186] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9191:9186] * PIXEL_SIZE && v_count < i_worm_y[9191:9186] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1532 < i_size && h_count >= i_worm_x[9197:9192] * PIXEL_SIZE && h_count < i_worm_x[9197:9192] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9197:9192] * PIXEL_SIZE && v_count < i_worm_y[9197:9192] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1533 < i_size && h_count >= i_worm_x[9203:9198] * PIXEL_SIZE && h_count < i_worm_x[9203:9198] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9203:9198] * PIXEL_SIZE && v_count < i_worm_y[9203:9198] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1534 < i_size && h_count >= i_worm_x[9209:9204] * PIXEL_SIZE && h_count < i_worm_x[9209:9204] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9209:9204] * PIXEL_SIZE && v_count < i_worm_y[9209:9204] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1535 < i_size && h_count >= i_worm_x[9215:9210] * PIXEL_SIZE && h_count < i_worm_x[9215:9210] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9215:9210] * PIXEL_SIZE && v_count < i_worm_y[9215:9210] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1536 < i_size && h_count >= i_worm_x[9221:9216] * PIXEL_SIZE && h_count < i_worm_x[9221:9216] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9221:9216] * PIXEL_SIZE && v_count < i_worm_y[9221:9216] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1537 < i_size && h_count >= i_worm_x[9227:9222] * PIXEL_SIZE && h_count < i_worm_x[9227:9222] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9227:9222] * PIXEL_SIZE && v_count < i_worm_y[9227:9222] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1538 < i_size && h_count >= i_worm_x[9233:9228] * PIXEL_SIZE && h_count < i_worm_x[9233:9228] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9233:9228] * PIXEL_SIZE && v_count < i_worm_y[9233:9228] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1539 < i_size && h_count >= i_worm_x[9239:9234] * PIXEL_SIZE && h_count < i_worm_x[9239:9234] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9239:9234] * PIXEL_SIZE && v_count < i_worm_y[9239:9234] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1540 < i_size && h_count >= i_worm_x[9245:9240] * PIXEL_SIZE && h_count < i_worm_x[9245:9240] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9245:9240] * PIXEL_SIZE && v_count < i_worm_y[9245:9240] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1541 < i_size && h_count >= i_worm_x[9251:9246] * PIXEL_SIZE && h_count < i_worm_x[9251:9246] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9251:9246] * PIXEL_SIZE && v_count < i_worm_y[9251:9246] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1542 < i_size && h_count >= i_worm_x[9257:9252] * PIXEL_SIZE && h_count < i_worm_x[9257:9252] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9257:9252] * PIXEL_SIZE && v_count < i_worm_y[9257:9252] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1543 < i_size && h_count >= i_worm_x[9263:9258] * PIXEL_SIZE && h_count < i_worm_x[9263:9258] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9263:9258] * PIXEL_SIZE && v_count < i_worm_y[9263:9258] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1544 < i_size && h_count >= i_worm_x[9269:9264] * PIXEL_SIZE && h_count < i_worm_x[9269:9264] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9269:9264] * PIXEL_SIZE && v_count < i_worm_y[9269:9264] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1545 < i_size && h_count >= i_worm_x[9275:9270] * PIXEL_SIZE && h_count < i_worm_x[9275:9270] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9275:9270] * PIXEL_SIZE && v_count < i_worm_y[9275:9270] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1546 < i_size && h_count >= i_worm_x[9281:9276] * PIXEL_SIZE && h_count < i_worm_x[9281:9276] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9281:9276] * PIXEL_SIZE && v_count < i_worm_y[9281:9276] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1547 < i_size && h_count >= i_worm_x[9287:9282] * PIXEL_SIZE && h_count < i_worm_x[9287:9282] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9287:9282] * PIXEL_SIZE && v_count < i_worm_y[9287:9282] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1548 < i_size && h_count >= i_worm_x[9293:9288] * PIXEL_SIZE && h_count < i_worm_x[9293:9288] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9293:9288] * PIXEL_SIZE && v_count < i_worm_y[9293:9288] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1549 < i_size && h_count >= i_worm_x[9299:9294] * PIXEL_SIZE && h_count < i_worm_x[9299:9294] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9299:9294] * PIXEL_SIZE && v_count < i_worm_y[9299:9294] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1550 < i_size && h_count >= i_worm_x[9305:9300] * PIXEL_SIZE && h_count < i_worm_x[9305:9300] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9305:9300] * PIXEL_SIZE && v_count < i_worm_y[9305:9300] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1551 < i_size && h_count >= i_worm_x[9311:9306] * PIXEL_SIZE && h_count < i_worm_x[9311:9306] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9311:9306] * PIXEL_SIZE && v_count < i_worm_y[9311:9306] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1552 < i_size && h_count >= i_worm_x[9317:9312] * PIXEL_SIZE && h_count < i_worm_x[9317:9312] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9317:9312] * PIXEL_SIZE && v_count < i_worm_y[9317:9312] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1553 < i_size && h_count >= i_worm_x[9323:9318] * PIXEL_SIZE && h_count < i_worm_x[9323:9318] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9323:9318] * PIXEL_SIZE && v_count < i_worm_y[9323:9318] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1554 < i_size && h_count >= i_worm_x[9329:9324] * PIXEL_SIZE && h_count < i_worm_x[9329:9324] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9329:9324] * PIXEL_SIZE && v_count < i_worm_y[9329:9324] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1555 < i_size && h_count >= i_worm_x[9335:9330] * PIXEL_SIZE && h_count < i_worm_x[9335:9330] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9335:9330] * PIXEL_SIZE && v_count < i_worm_y[9335:9330] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1556 < i_size && h_count >= i_worm_x[9341:9336] * PIXEL_SIZE && h_count < i_worm_x[9341:9336] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9341:9336] * PIXEL_SIZE && v_count < i_worm_y[9341:9336] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1557 < i_size && h_count >= i_worm_x[9347:9342] * PIXEL_SIZE && h_count < i_worm_x[9347:9342] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9347:9342] * PIXEL_SIZE && v_count < i_worm_y[9347:9342] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1558 < i_size && h_count >= i_worm_x[9353:9348] * PIXEL_SIZE && h_count < i_worm_x[9353:9348] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9353:9348] * PIXEL_SIZE && v_count < i_worm_y[9353:9348] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1559 < i_size && h_count >= i_worm_x[9359:9354] * PIXEL_SIZE && h_count < i_worm_x[9359:9354] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9359:9354] * PIXEL_SIZE && v_count < i_worm_y[9359:9354] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1560 < i_size && h_count >= i_worm_x[9365:9360] * PIXEL_SIZE && h_count < i_worm_x[9365:9360] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9365:9360] * PIXEL_SIZE && v_count < i_worm_y[9365:9360] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1561 < i_size && h_count >= i_worm_x[9371:9366] * PIXEL_SIZE && h_count < i_worm_x[9371:9366] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9371:9366] * PIXEL_SIZE && v_count < i_worm_y[9371:9366] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1562 < i_size && h_count >= i_worm_x[9377:9372] * PIXEL_SIZE && h_count < i_worm_x[9377:9372] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9377:9372] * PIXEL_SIZE && v_count < i_worm_y[9377:9372] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1563 < i_size && h_count >= i_worm_x[9383:9378] * PIXEL_SIZE && h_count < i_worm_x[9383:9378] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9383:9378] * PIXEL_SIZE && v_count < i_worm_y[9383:9378] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1564 < i_size && h_count >= i_worm_x[9389:9384] * PIXEL_SIZE && h_count < i_worm_x[9389:9384] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9389:9384] * PIXEL_SIZE && v_count < i_worm_y[9389:9384] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1565 < i_size && h_count >= i_worm_x[9395:9390] * PIXEL_SIZE && h_count < i_worm_x[9395:9390] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9395:9390] * PIXEL_SIZE && v_count < i_worm_y[9395:9390] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1566 < i_size && h_count >= i_worm_x[9401:9396] * PIXEL_SIZE && h_count < i_worm_x[9401:9396] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9401:9396] * PIXEL_SIZE && v_count < i_worm_y[9401:9396] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1567 < i_size && h_count >= i_worm_x[9407:9402] * PIXEL_SIZE && h_count < i_worm_x[9407:9402] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9407:9402] * PIXEL_SIZE && v_count < i_worm_y[9407:9402] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1568 < i_size && h_count >= i_worm_x[9413:9408] * PIXEL_SIZE && h_count < i_worm_x[9413:9408] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9413:9408] * PIXEL_SIZE && v_count < i_worm_y[9413:9408] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1569 < i_size && h_count >= i_worm_x[9419:9414] * PIXEL_SIZE && h_count < i_worm_x[9419:9414] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9419:9414] * PIXEL_SIZE && v_count < i_worm_y[9419:9414] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1570 < i_size && h_count >= i_worm_x[9425:9420] * PIXEL_SIZE && h_count < i_worm_x[9425:9420] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9425:9420] * PIXEL_SIZE && v_count < i_worm_y[9425:9420] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1571 < i_size && h_count >= i_worm_x[9431:9426] * PIXEL_SIZE && h_count < i_worm_x[9431:9426] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9431:9426] * PIXEL_SIZE && v_count < i_worm_y[9431:9426] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1572 < i_size && h_count >= i_worm_x[9437:9432] * PIXEL_SIZE && h_count < i_worm_x[9437:9432] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9437:9432] * PIXEL_SIZE && v_count < i_worm_y[9437:9432] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1573 < i_size && h_count >= i_worm_x[9443:9438] * PIXEL_SIZE && h_count < i_worm_x[9443:9438] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9443:9438] * PIXEL_SIZE && v_count < i_worm_y[9443:9438] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1574 < i_size && h_count >= i_worm_x[9449:9444] * PIXEL_SIZE && h_count < i_worm_x[9449:9444] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9449:9444] * PIXEL_SIZE && v_count < i_worm_y[9449:9444] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1575 < i_size && h_count >= i_worm_x[9455:9450] * PIXEL_SIZE && h_count < i_worm_x[9455:9450] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9455:9450] * PIXEL_SIZE && v_count < i_worm_y[9455:9450] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1576 < i_size && h_count >= i_worm_x[9461:9456] * PIXEL_SIZE && h_count < i_worm_x[9461:9456] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9461:9456] * PIXEL_SIZE && v_count < i_worm_y[9461:9456] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1577 < i_size && h_count >= i_worm_x[9467:9462] * PIXEL_SIZE && h_count < i_worm_x[9467:9462] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9467:9462] * PIXEL_SIZE && v_count < i_worm_y[9467:9462] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1578 < i_size && h_count >= i_worm_x[9473:9468] * PIXEL_SIZE && h_count < i_worm_x[9473:9468] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9473:9468] * PIXEL_SIZE && v_count < i_worm_y[9473:9468] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1579 < i_size && h_count >= i_worm_x[9479:9474] * PIXEL_SIZE && h_count < i_worm_x[9479:9474] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9479:9474] * PIXEL_SIZE && v_count < i_worm_y[9479:9474] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1580 < i_size && h_count >= i_worm_x[9485:9480] * PIXEL_SIZE && h_count < i_worm_x[9485:9480] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9485:9480] * PIXEL_SIZE && v_count < i_worm_y[9485:9480] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1581 < i_size && h_count >= i_worm_x[9491:9486] * PIXEL_SIZE && h_count < i_worm_x[9491:9486] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9491:9486] * PIXEL_SIZE && v_count < i_worm_y[9491:9486] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1582 < i_size && h_count >= i_worm_x[9497:9492] * PIXEL_SIZE && h_count < i_worm_x[9497:9492] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9497:9492] * PIXEL_SIZE && v_count < i_worm_y[9497:9492] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1583 < i_size && h_count >= i_worm_x[9503:9498] * PIXEL_SIZE && h_count < i_worm_x[9503:9498] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9503:9498] * PIXEL_SIZE && v_count < i_worm_y[9503:9498] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1584 < i_size && h_count >= i_worm_x[9509:9504] * PIXEL_SIZE && h_count < i_worm_x[9509:9504] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9509:9504] * PIXEL_SIZE && v_count < i_worm_y[9509:9504] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1585 < i_size && h_count >= i_worm_x[9515:9510] * PIXEL_SIZE && h_count < i_worm_x[9515:9510] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9515:9510] * PIXEL_SIZE && v_count < i_worm_y[9515:9510] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1586 < i_size && h_count >= i_worm_x[9521:9516] * PIXEL_SIZE && h_count < i_worm_x[9521:9516] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9521:9516] * PIXEL_SIZE && v_count < i_worm_y[9521:9516] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1587 < i_size && h_count >= i_worm_x[9527:9522] * PIXEL_SIZE && h_count < i_worm_x[9527:9522] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9527:9522] * PIXEL_SIZE && v_count < i_worm_y[9527:9522] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1588 < i_size && h_count >= i_worm_x[9533:9528] * PIXEL_SIZE && h_count < i_worm_x[9533:9528] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9533:9528] * PIXEL_SIZE && v_count < i_worm_y[9533:9528] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1589 < i_size && h_count >= i_worm_x[9539:9534] * PIXEL_SIZE && h_count < i_worm_x[9539:9534] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9539:9534] * PIXEL_SIZE && v_count < i_worm_y[9539:9534] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1590 < i_size && h_count >= i_worm_x[9545:9540] * PIXEL_SIZE && h_count < i_worm_x[9545:9540] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9545:9540] * PIXEL_SIZE && v_count < i_worm_y[9545:9540] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1591 < i_size && h_count >= i_worm_x[9551:9546] * PIXEL_SIZE && h_count < i_worm_x[9551:9546] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9551:9546] * PIXEL_SIZE && v_count < i_worm_y[9551:9546] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1592 < i_size && h_count >= i_worm_x[9557:9552] * PIXEL_SIZE && h_count < i_worm_x[9557:9552] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9557:9552] * PIXEL_SIZE && v_count < i_worm_y[9557:9552] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1593 < i_size && h_count >= i_worm_x[9563:9558] * PIXEL_SIZE && h_count < i_worm_x[9563:9558] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9563:9558] * PIXEL_SIZE && v_count < i_worm_y[9563:9558] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1594 < i_size && h_count >= i_worm_x[9569:9564] * PIXEL_SIZE && h_count < i_worm_x[9569:9564] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9569:9564] * PIXEL_SIZE && v_count < i_worm_y[9569:9564] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1595 < i_size && h_count >= i_worm_x[9575:9570] * PIXEL_SIZE && h_count < i_worm_x[9575:9570] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9575:9570] * PIXEL_SIZE && v_count < i_worm_y[9575:9570] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1596 < i_size && h_count >= i_worm_x[9581:9576] * PIXEL_SIZE && h_count < i_worm_x[9581:9576] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9581:9576] * PIXEL_SIZE && v_count < i_worm_y[9581:9576] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1597 < i_size && h_count >= i_worm_x[9587:9582] * PIXEL_SIZE && h_count < i_worm_x[9587:9582] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9587:9582] * PIXEL_SIZE && v_count < i_worm_y[9587:9582] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1598 < i_size && h_count >= i_worm_x[9593:9588] * PIXEL_SIZE && h_count < i_worm_x[9593:9588] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9593:9588] * PIXEL_SIZE && v_count < i_worm_y[9593:9588] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1599 < i_size && h_count >= i_worm_x[9599:9594] * PIXEL_SIZE && h_count < i_worm_x[9599:9594] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9599:9594] * PIXEL_SIZE && v_count < i_worm_y[9599:9594] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1600 < i_size && h_count >= i_worm_x[9605:9600] * PIXEL_SIZE && h_count < i_worm_x[9605:9600] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9605:9600] * PIXEL_SIZE && v_count < i_worm_y[9605:9600] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1601 < i_size && h_count >= i_worm_x[9611:9606] * PIXEL_SIZE && h_count < i_worm_x[9611:9606] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9611:9606] * PIXEL_SIZE && v_count < i_worm_y[9611:9606] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1602 < i_size && h_count >= i_worm_x[9617:9612] * PIXEL_SIZE && h_count < i_worm_x[9617:9612] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9617:9612] * PIXEL_SIZE && v_count < i_worm_y[9617:9612] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1603 < i_size && h_count >= i_worm_x[9623:9618] * PIXEL_SIZE && h_count < i_worm_x[9623:9618] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9623:9618] * PIXEL_SIZE && v_count < i_worm_y[9623:9618] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1604 < i_size && h_count >= i_worm_x[9629:9624] * PIXEL_SIZE && h_count < i_worm_x[9629:9624] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9629:9624] * PIXEL_SIZE && v_count < i_worm_y[9629:9624] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1605 < i_size && h_count >= i_worm_x[9635:9630] * PIXEL_SIZE && h_count < i_worm_x[9635:9630] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9635:9630] * PIXEL_SIZE && v_count < i_worm_y[9635:9630] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1606 < i_size && h_count >= i_worm_x[9641:9636] * PIXEL_SIZE && h_count < i_worm_x[9641:9636] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9641:9636] * PIXEL_SIZE && v_count < i_worm_y[9641:9636] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1607 < i_size && h_count >= i_worm_x[9647:9642] * PIXEL_SIZE && h_count < i_worm_x[9647:9642] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9647:9642] * PIXEL_SIZE && v_count < i_worm_y[9647:9642] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1608 < i_size && h_count >= i_worm_x[9653:9648] * PIXEL_SIZE && h_count < i_worm_x[9653:9648] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9653:9648] * PIXEL_SIZE && v_count < i_worm_y[9653:9648] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1609 < i_size && h_count >= i_worm_x[9659:9654] * PIXEL_SIZE && h_count < i_worm_x[9659:9654] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9659:9654] * PIXEL_SIZE && v_count < i_worm_y[9659:9654] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1610 < i_size && h_count >= i_worm_x[9665:9660] * PIXEL_SIZE && h_count < i_worm_x[9665:9660] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9665:9660] * PIXEL_SIZE && v_count < i_worm_y[9665:9660] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1611 < i_size && h_count >= i_worm_x[9671:9666] * PIXEL_SIZE && h_count < i_worm_x[9671:9666] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9671:9666] * PIXEL_SIZE && v_count < i_worm_y[9671:9666] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1612 < i_size && h_count >= i_worm_x[9677:9672] * PIXEL_SIZE && h_count < i_worm_x[9677:9672] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9677:9672] * PIXEL_SIZE && v_count < i_worm_y[9677:9672] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1613 < i_size && h_count >= i_worm_x[9683:9678] * PIXEL_SIZE && h_count < i_worm_x[9683:9678] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9683:9678] * PIXEL_SIZE && v_count < i_worm_y[9683:9678] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1614 < i_size && h_count >= i_worm_x[9689:9684] * PIXEL_SIZE && h_count < i_worm_x[9689:9684] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9689:9684] * PIXEL_SIZE && v_count < i_worm_y[9689:9684] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1615 < i_size && h_count >= i_worm_x[9695:9690] * PIXEL_SIZE && h_count < i_worm_x[9695:9690] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9695:9690] * PIXEL_SIZE && v_count < i_worm_y[9695:9690] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1616 < i_size && h_count >= i_worm_x[9701:9696] * PIXEL_SIZE && h_count < i_worm_x[9701:9696] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9701:9696] * PIXEL_SIZE && v_count < i_worm_y[9701:9696] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1617 < i_size && h_count >= i_worm_x[9707:9702] * PIXEL_SIZE && h_count < i_worm_x[9707:9702] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9707:9702] * PIXEL_SIZE && v_count < i_worm_y[9707:9702] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1618 < i_size && h_count >= i_worm_x[9713:9708] * PIXEL_SIZE && h_count < i_worm_x[9713:9708] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9713:9708] * PIXEL_SIZE && v_count < i_worm_y[9713:9708] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1619 < i_size && h_count >= i_worm_x[9719:9714] * PIXEL_SIZE && h_count < i_worm_x[9719:9714] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9719:9714] * PIXEL_SIZE && v_count < i_worm_y[9719:9714] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1620 < i_size && h_count >= i_worm_x[9725:9720] * PIXEL_SIZE && h_count < i_worm_x[9725:9720] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9725:9720] * PIXEL_SIZE && v_count < i_worm_y[9725:9720] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1621 < i_size && h_count >= i_worm_x[9731:9726] * PIXEL_SIZE && h_count < i_worm_x[9731:9726] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9731:9726] * PIXEL_SIZE && v_count < i_worm_y[9731:9726] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1622 < i_size && h_count >= i_worm_x[9737:9732] * PIXEL_SIZE && h_count < i_worm_x[9737:9732] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9737:9732] * PIXEL_SIZE && v_count < i_worm_y[9737:9732] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1623 < i_size && h_count >= i_worm_x[9743:9738] * PIXEL_SIZE && h_count < i_worm_x[9743:9738] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9743:9738] * PIXEL_SIZE && v_count < i_worm_y[9743:9738] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1624 < i_size && h_count >= i_worm_x[9749:9744] * PIXEL_SIZE && h_count < i_worm_x[9749:9744] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9749:9744] * PIXEL_SIZE && v_count < i_worm_y[9749:9744] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1625 < i_size && h_count >= i_worm_x[9755:9750] * PIXEL_SIZE && h_count < i_worm_x[9755:9750] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9755:9750] * PIXEL_SIZE && v_count < i_worm_y[9755:9750] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1626 < i_size && h_count >= i_worm_x[9761:9756] * PIXEL_SIZE && h_count < i_worm_x[9761:9756] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9761:9756] * PIXEL_SIZE && v_count < i_worm_y[9761:9756] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1627 < i_size && h_count >= i_worm_x[9767:9762] * PIXEL_SIZE && h_count < i_worm_x[9767:9762] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9767:9762] * PIXEL_SIZE && v_count < i_worm_y[9767:9762] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1628 < i_size && h_count >= i_worm_x[9773:9768] * PIXEL_SIZE && h_count < i_worm_x[9773:9768] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9773:9768] * PIXEL_SIZE && v_count < i_worm_y[9773:9768] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1629 < i_size && h_count >= i_worm_x[9779:9774] * PIXEL_SIZE && h_count < i_worm_x[9779:9774] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9779:9774] * PIXEL_SIZE && v_count < i_worm_y[9779:9774] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1630 < i_size && h_count >= i_worm_x[9785:9780] * PIXEL_SIZE && h_count < i_worm_x[9785:9780] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9785:9780] * PIXEL_SIZE && v_count < i_worm_y[9785:9780] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1631 < i_size && h_count >= i_worm_x[9791:9786] * PIXEL_SIZE && h_count < i_worm_x[9791:9786] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9791:9786] * PIXEL_SIZE && v_count < i_worm_y[9791:9786] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1632 < i_size && h_count >= i_worm_x[9797:9792] * PIXEL_SIZE && h_count < i_worm_x[9797:9792] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9797:9792] * PIXEL_SIZE && v_count < i_worm_y[9797:9792] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1633 < i_size && h_count >= i_worm_x[9803:9798] * PIXEL_SIZE && h_count < i_worm_x[9803:9798] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9803:9798] * PIXEL_SIZE && v_count < i_worm_y[9803:9798] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1634 < i_size && h_count >= i_worm_x[9809:9804] * PIXEL_SIZE && h_count < i_worm_x[9809:9804] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9809:9804] * PIXEL_SIZE && v_count < i_worm_y[9809:9804] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1635 < i_size && h_count >= i_worm_x[9815:9810] * PIXEL_SIZE && h_count < i_worm_x[9815:9810] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9815:9810] * PIXEL_SIZE && v_count < i_worm_y[9815:9810] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1636 < i_size && h_count >= i_worm_x[9821:9816] * PIXEL_SIZE && h_count < i_worm_x[9821:9816] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9821:9816] * PIXEL_SIZE && v_count < i_worm_y[9821:9816] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1637 < i_size && h_count >= i_worm_x[9827:9822] * PIXEL_SIZE && h_count < i_worm_x[9827:9822] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9827:9822] * PIXEL_SIZE && v_count < i_worm_y[9827:9822] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1638 < i_size && h_count >= i_worm_x[9833:9828] * PIXEL_SIZE && h_count < i_worm_x[9833:9828] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9833:9828] * PIXEL_SIZE && v_count < i_worm_y[9833:9828] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1639 < i_size && h_count >= i_worm_x[9839:9834] * PIXEL_SIZE && h_count < i_worm_x[9839:9834] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9839:9834] * PIXEL_SIZE && v_count < i_worm_y[9839:9834] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1640 < i_size && h_count >= i_worm_x[9845:9840] * PIXEL_SIZE && h_count < i_worm_x[9845:9840] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9845:9840] * PIXEL_SIZE && v_count < i_worm_y[9845:9840] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1641 < i_size && h_count >= i_worm_x[9851:9846] * PIXEL_SIZE && h_count < i_worm_x[9851:9846] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9851:9846] * PIXEL_SIZE && v_count < i_worm_y[9851:9846] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1642 < i_size && h_count >= i_worm_x[9857:9852] * PIXEL_SIZE && h_count < i_worm_x[9857:9852] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9857:9852] * PIXEL_SIZE && v_count < i_worm_y[9857:9852] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1643 < i_size && h_count >= i_worm_x[9863:9858] * PIXEL_SIZE && h_count < i_worm_x[9863:9858] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9863:9858] * PIXEL_SIZE && v_count < i_worm_y[9863:9858] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1644 < i_size && h_count >= i_worm_x[9869:9864] * PIXEL_SIZE && h_count < i_worm_x[9869:9864] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9869:9864] * PIXEL_SIZE && v_count < i_worm_y[9869:9864] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1645 < i_size && h_count >= i_worm_x[9875:9870] * PIXEL_SIZE && h_count < i_worm_x[9875:9870] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9875:9870] * PIXEL_SIZE && v_count < i_worm_y[9875:9870] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1646 < i_size && h_count >= i_worm_x[9881:9876] * PIXEL_SIZE && h_count < i_worm_x[9881:9876] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9881:9876] * PIXEL_SIZE && v_count < i_worm_y[9881:9876] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1647 < i_size && h_count >= i_worm_x[9887:9882] * PIXEL_SIZE && h_count < i_worm_x[9887:9882] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9887:9882] * PIXEL_SIZE && v_count < i_worm_y[9887:9882] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1648 < i_size && h_count >= i_worm_x[9893:9888] * PIXEL_SIZE && h_count < i_worm_x[9893:9888] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9893:9888] * PIXEL_SIZE && v_count < i_worm_y[9893:9888] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1649 < i_size && h_count >= i_worm_x[9899:9894] * PIXEL_SIZE && h_count < i_worm_x[9899:9894] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9899:9894] * PIXEL_SIZE && v_count < i_worm_y[9899:9894] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1650 < i_size && h_count >= i_worm_x[9905:9900] * PIXEL_SIZE && h_count < i_worm_x[9905:9900] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9905:9900] * PIXEL_SIZE && v_count < i_worm_y[9905:9900] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1651 < i_size && h_count >= i_worm_x[9911:9906] * PIXEL_SIZE && h_count < i_worm_x[9911:9906] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9911:9906] * PIXEL_SIZE && v_count < i_worm_y[9911:9906] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1652 < i_size && h_count >= i_worm_x[9917:9912] * PIXEL_SIZE && h_count < i_worm_x[9917:9912] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9917:9912] * PIXEL_SIZE && v_count < i_worm_y[9917:9912] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1653 < i_size && h_count >= i_worm_x[9923:9918] * PIXEL_SIZE && h_count < i_worm_x[9923:9918] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9923:9918] * PIXEL_SIZE && v_count < i_worm_y[9923:9918] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1654 < i_size && h_count >= i_worm_x[9929:9924] * PIXEL_SIZE && h_count < i_worm_x[9929:9924] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9929:9924] * PIXEL_SIZE && v_count < i_worm_y[9929:9924] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1655 < i_size && h_count >= i_worm_x[9935:9930] * PIXEL_SIZE && h_count < i_worm_x[9935:9930] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9935:9930] * PIXEL_SIZE && v_count < i_worm_y[9935:9930] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1656 < i_size && h_count >= i_worm_x[9941:9936] * PIXEL_SIZE && h_count < i_worm_x[9941:9936] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9941:9936] * PIXEL_SIZE && v_count < i_worm_y[9941:9936] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1657 < i_size && h_count >= i_worm_x[9947:9942] * PIXEL_SIZE && h_count < i_worm_x[9947:9942] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9947:9942] * PIXEL_SIZE && v_count < i_worm_y[9947:9942] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1658 < i_size && h_count >= i_worm_x[9953:9948] * PIXEL_SIZE && h_count < i_worm_x[9953:9948] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9953:9948] * PIXEL_SIZE && v_count < i_worm_y[9953:9948] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1659 < i_size && h_count >= i_worm_x[9959:9954] * PIXEL_SIZE && h_count < i_worm_x[9959:9954] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9959:9954] * PIXEL_SIZE && v_count < i_worm_y[9959:9954] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1660 < i_size && h_count >= i_worm_x[9965:9960] * PIXEL_SIZE && h_count < i_worm_x[9965:9960] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9965:9960] * PIXEL_SIZE && v_count < i_worm_y[9965:9960] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1661 < i_size && h_count >= i_worm_x[9971:9966] * PIXEL_SIZE && h_count < i_worm_x[9971:9966] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9971:9966] * PIXEL_SIZE && v_count < i_worm_y[9971:9966] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1662 < i_size && h_count >= i_worm_x[9977:9972] * PIXEL_SIZE && h_count < i_worm_x[9977:9972] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9977:9972] * PIXEL_SIZE && v_count < i_worm_y[9977:9972] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1663 < i_size && h_count >= i_worm_x[9983:9978] * PIXEL_SIZE && h_count < i_worm_x[9983:9978] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9983:9978] * PIXEL_SIZE && v_count < i_worm_y[9983:9978] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1664 < i_size && h_count >= i_worm_x[9989:9984] * PIXEL_SIZE && h_count < i_worm_x[9989:9984] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9989:9984] * PIXEL_SIZE && v_count < i_worm_y[9989:9984] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1665 < i_size && h_count >= i_worm_x[9995:9990] * PIXEL_SIZE && h_count < i_worm_x[9995:9990] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[9995:9990] * PIXEL_SIZE && v_count < i_worm_y[9995:9990] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1666 < i_size && h_count >= i_worm_x[10001:9996] * PIXEL_SIZE && h_count < i_worm_x[10001:9996] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10001:9996] * PIXEL_SIZE && v_count < i_worm_y[10001:9996] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1667 < i_size && h_count >= i_worm_x[10007:10002] * PIXEL_SIZE && h_count < i_worm_x[10007:10002] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10007:10002] * PIXEL_SIZE && v_count < i_worm_y[10007:10002] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1668 < i_size && h_count >= i_worm_x[10013:10008] * PIXEL_SIZE && h_count < i_worm_x[10013:10008] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10013:10008] * PIXEL_SIZE && v_count < i_worm_y[10013:10008] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1669 < i_size && h_count >= i_worm_x[10019:10014] * PIXEL_SIZE && h_count < i_worm_x[10019:10014] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10019:10014] * PIXEL_SIZE && v_count < i_worm_y[10019:10014] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1670 < i_size && h_count >= i_worm_x[10025:10020] * PIXEL_SIZE && h_count < i_worm_x[10025:10020] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10025:10020] * PIXEL_SIZE && v_count < i_worm_y[10025:10020] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1671 < i_size && h_count >= i_worm_x[10031:10026] * PIXEL_SIZE && h_count < i_worm_x[10031:10026] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10031:10026] * PIXEL_SIZE && v_count < i_worm_y[10031:10026] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1672 < i_size && h_count >= i_worm_x[10037:10032] * PIXEL_SIZE && h_count < i_worm_x[10037:10032] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10037:10032] * PIXEL_SIZE && v_count < i_worm_y[10037:10032] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1673 < i_size && h_count >= i_worm_x[10043:10038] * PIXEL_SIZE && h_count < i_worm_x[10043:10038] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10043:10038] * PIXEL_SIZE && v_count < i_worm_y[10043:10038] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1674 < i_size && h_count >= i_worm_x[10049:10044] * PIXEL_SIZE && h_count < i_worm_x[10049:10044] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10049:10044] * PIXEL_SIZE && v_count < i_worm_y[10049:10044] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1675 < i_size && h_count >= i_worm_x[10055:10050] * PIXEL_SIZE && h_count < i_worm_x[10055:10050] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10055:10050] * PIXEL_SIZE && v_count < i_worm_y[10055:10050] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1676 < i_size && h_count >= i_worm_x[10061:10056] * PIXEL_SIZE && h_count < i_worm_x[10061:10056] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10061:10056] * PIXEL_SIZE && v_count < i_worm_y[10061:10056] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1677 < i_size && h_count >= i_worm_x[10067:10062] * PIXEL_SIZE && h_count < i_worm_x[10067:10062] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10067:10062] * PIXEL_SIZE && v_count < i_worm_y[10067:10062] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1678 < i_size && h_count >= i_worm_x[10073:10068] * PIXEL_SIZE && h_count < i_worm_x[10073:10068] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10073:10068] * PIXEL_SIZE && v_count < i_worm_y[10073:10068] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1679 < i_size && h_count >= i_worm_x[10079:10074] * PIXEL_SIZE && h_count < i_worm_x[10079:10074] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10079:10074] * PIXEL_SIZE && v_count < i_worm_y[10079:10074] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1680 < i_size && h_count >= i_worm_x[10085:10080] * PIXEL_SIZE && h_count < i_worm_x[10085:10080] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10085:10080] * PIXEL_SIZE && v_count < i_worm_y[10085:10080] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1681 < i_size && h_count >= i_worm_x[10091:10086] * PIXEL_SIZE && h_count < i_worm_x[10091:10086] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10091:10086] * PIXEL_SIZE && v_count < i_worm_y[10091:10086] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1682 < i_size && h_count >= i_worm_x[10097:10092] * PIXEL_SIZE && h_count < i_worm_x[10097:10092] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10097:10092] * PIXEL_SIZE && v_count < i_worm_y[10097:10092] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1683 < i_size && h_count >= i_worm_x[10103:10098] * PIXEL_SIZE && h_count < i_worm_x[10103:10098] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10103:10098] * PIXEL_SIZE && v_count < i_worm_y[10103:10098] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1684 < i_size && h_count >= i_worm_x[10109:10104] * PIXEL_SIZE && h_count < i_worm_x[10109:10104] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10109:10104] * PIXEL_SIZE && v_count < i_worm_y[10109:10104] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1685 < i_size && h_count >= i_worm_x[10115:10110] * PIXEL_SIZE && h_count < i_worm_x[10115:10110] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10115:10110] * PIXEL_SIZE && v_count < i_worm_y[10115:10110] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1686 < i_size && h_count >= i_worm_x[10121:10116] * PIXEL_SIZE && h_count < i_worm_x[10121:10116] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10121:10116] * PIXEL_SIZE && v_count < i_worm_y[10121:10116] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1687 < i_size && h_count >= i_worm_x[10127:10122] * PIXEL_SIZE && h_count < i_worm_x[10127:10122] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10127:10122] * PIXEL_SIZE && v_count < i_worm_y[10127:10122] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1688 < i_size && h_count >= i_worm_x[10133:10128] * PIXEL_SIZE && h_count < i_worm_x[10133:10128] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10133:10128] * PIXEL_SIZE && v_count < i_worm_y[10133:10128] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1689 < i_size && h_count >= i_worm_x[10139:10134] * PIXEL_SIZE && h_count < i_worm_x[10139:10134] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10139:10134] * PIXEL_SIZE && v_count < i_worm_y[10139:10134] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1690 < i_size && h_count >= i_worm_x[10145:10140] * PIXEL_SIZE && h_count < i_worm_x[10145:10140] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10145:10140] * PIXEL_SIZE && v_count < i_worm_y[10145:10140] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1691 < i_size && h_count >= i_worm_x[10151:10146] * PIXEL_SIZE && h_count < i_worm_x[10151:10146] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10151:10146] * PIXEL_SIZE && v_count < i_worm_y[10151:10146] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1692 < i_size && h_count >= i_worm_x[10157:10152] * PIXEL_SIZE && h_count < i_worm_x[10157:10152] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10157:10152] * PIXEL_SIZE && v_count < i_worm_y[10157:10152] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1693 < i_size && h_count >= i_worm_x[10163:10158] * PIXEL_SIZE && h_count < i_worm_x[10163:10158] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10163:10158] * PIXEL_SIZE && v_count < i_worm_y[10163:10158] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1694 < i_size && h_count >= i_worm_x[10169:10164] * PIXEL_SIZE && h_count < i_worm_x[10169:10164] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10169:10164] * PIXEL_SIZE && v_count < i_worm_y[10169:10164] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1695 < i_size && h_count >= i_worm_x[10175:10170] * PIXEL_SIZE && h_count < i_worm_x[10175:10170] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10175:10170] * PIXEL_SIZE && v_count < i_worm_y[10175:10170] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1696 < i_size && h_count >= i_worm_x[10181:10176] * PIXEL_SIZE && h_count < i_worm_x[10181:10176] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10181:10176] * PIXEL_SIZE && v_count < i_worm_y[10181:10176] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1697 < i_size && h_count >= i_worm_x[10187:10182] * PIXEL_SIZE && h_count < i_worm_x[10187:10182] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10187:10182] * PIXEL_SIZE && v_count < i_worm_y[10187:10182] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1698 < i_size && h_count >= i_worm_x[10193:10188] * PIXEL_SIZE && h_count < i_worm_x[10193:10188] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10193:10188] * PIXEL_SIZE && v_count < i_worm_y[10193:10188] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1699 < i_size && h_count >= i_worm_x[10199:10194] * PIXEL_SIZE && h_count < i_worm_x[10199:10194] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10199:10194] * PIXEL_SIZE && v_count < i_worm_y[10199:10194] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1700 < i_size && h_count >= i_worm_x[10205:10200] * PIXEL_SIZE && h_count < i_worm_x[10205:10200] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10205:10200] * PIXEL_SIZE && v_count < i_worm_y[10205:10200] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1701 < i_size && h_count >= i_worm_x[10211:10206] * PIXEL_SIZE && h_count < i_worm_x[10211:10206] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10211:10206] * PIXEL_SIZE && v_count < i_worm_y[10211:10206] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1702 < i_size && h_count >= i_worm_x[10217:10212] * PIXEL_SIZE && h_count < i_worm_x[10217:10212] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10217:10212] * PIXEL_SIZE && v_count < i_worm_y[10217:10212] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1703 < i_size && h_count >= i_worm_x[10223:10218] * PIXEL_SIZE && h_count < i_worm_x[10223:10218] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10223:10218] * PIXEL_SIZE && v_count < i_worm_y[10223:10218] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1704 < i_size && h_count >= i_worm_x[10229:10224] * PIXEL_SIZE && h_count < i_worm_x[10229:10224] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10229:10224] * PIXEL_SIZE && v_count < i_worm_y[10229:10224] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1705 < i_size && h_count >= i_worm_x[10235:10230] * PIXEL_SIZE && h_count < i_worm_x[10235:10230] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10235:10230] * PIXEL_SIZE && v_count < i_worm_y[10235:10230] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1706 < i_size && h_count >= i_worm_x[10241:10236] * PIXEL_SIZE && h_count < i_worm_x[10241:10236] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10241:10236] * PIXEL_SIZE && v_count < i_worm_y[10241:10236] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1707 < i_size && h_count >= i_worm_x[10247:10242] * PIXEL_SIZE && h_count < i_worm_x[10247:10242] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10247:10242] * PIXEL_SIZE && v_count < i_worm_y[10247:10242] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1708 < i_size && h_count >= i_worm_x[10253:10248] * PIXEL_SIZE && h_count < i_worm_x[10253:10248] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10253:10248] * PIXEL_SIZE && v_count < i_worm_y[10253:10248] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1709 < i_size && h_count >= i_worm_x[10259:10254] * PIXEL_SIZE && h_count < i_worm_x[10259:10254] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10259:10254] * PIXEL_SIZE && v_count < i_worm_y[10259:10254] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1710 < i_size && h_count >= i_worm_x[10265:10260] * PIXEL_SIZE && h_count < i_worm_x[10265:10260] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10265:10260] * PIXEL_SIZE && v_count < i_worm_y[10265:10260] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1711 < i_size && h_count >= i_worm_x[10271:10266] * PIXEL_SIZE && h_count < i_worm_x[10271:10266] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10271:10266] * PIXEL_SIZE && v_count < i_worm_y[10271:10266] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1712 < i_size && h_count >= i_worm_x[10277:10272] * PIXEL_SIZE && h_count < i_worm_x[10277:10272] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10277:10272] * PIXEL_SIZE && v_count < i_worm_y[10277:10272] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1713 < i_size && h_count >= i_worm_x[10283:10278] * PIXEL_SIZE && h_count < i_worm_x[10283:10278] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10283:10278] * PIXEL_SIZE && v_count < i_worm_y[10283:10278] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1714 < i_size && h_count >= i_worm_x[10289:10284] * PIXEL_SIZE && h_count < i_worm_x[10289:10284] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10289:10284] * PIXEL_SIZE && v_count < i_worm_y[10289:10284] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1715 < i_size && h_count >= i_worm_x[10295:10290] * PIXEL_SIZE && h_count < i_worm_x[10295:10290] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10295:10290] * PIXEL_SIZE && v_count < i_worm_y[10295:10290] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1716 < i_size && h_count >= i_worm_x[10301:10296] * PIXEL_SIZE && h_count < i_worm_x[10301:10296] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10301:10296] * PIXEL_SIZE && v_count < i_worm_y[10301:10296] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1717 < i_size && h_count >= i_worm_x[10307:10302] * PIXEL_SIZE && h_count < i_worm_x[10307:10302] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10307:10302] * PIXEL_SIZE && v_count < i_worm_y[10307:10302] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1718 < i_size && h_count >= i_worm_x[10313:10308] * PIXEL_SIZE && h_count < i_worm_x[10313:10308] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10313:10308] * PIXEL_SIZE && v_count < i_worm_y[10313:10308] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1719 < i_size && h_count >= i_worm_x[10319:10314] * PIXEL_SIZE && h_count < i_worm_x[10319:10314] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10319:10314] * PIXEL_SIZE && v_count < i_worm_y[10319:10314] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1720 < i_size && h_count >= i_worm_x[10325:10320] * PIXEL_SIZE && h_count < i_worm_x[10325:10320] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10325:10320] * PIXEL_SIZE && v_count < i_worm_y[10325:10320] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1721 < i_size && h_count >= i_worm_x[10331:10326] * PIXEL_SIZE && h_count < i_worm_x[10331:10326] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10331:10326] * PIXEL_SIZE && v_count < i_worm_y[10331:10326] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1722 < i_size && h_count >= i_worm_x[10337:10332] * PIXEL_SIZE && h_count < i_worm_x[10337:10332] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10337:10332] * PIXEL_SIZE && v_count < i_worm_y[10337:10332] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1723 < i_size && h_count >= i_worm_x[10343:10338] * PIXEL_SIZE && h_count < i_worm_x[10343:10338] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10343:10338] * PIXEL_SIZE && v_count < i_worm_y[10343:10338] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1724 < i_size && h_count >= i_worm_x[10349:10344] * PIXEL_SIZE && h_count < i_worm_x[10349:10344] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10349:10344] * PIXEL_SIZE && v_count < i_worm_y[10349:10344] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1725 < i_size && h_count >= i_worm_x[10355:10350] * PIXEL_SIZE && h_count < i_worm_x[10355:10350] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10355:10350] * PIXEL_SIZE && v_count < i_worm_y[10355:10350] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1726 < i_size && h_count >= i_worm_x[10361:10356] * PIXEL_SIZE && h_count < i_worm_x[10361:10356] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10361:10356] * PIXEL_SIZE && v_count < i_worm_y[10361:10356] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1727 < i_size && h_count >= i_worm_x[10367:10362] * PIXEL_SIZE && h_count < i_worm_x[10367:10362] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10367:10362] * PIXEL_SIZE && v_count < i_worm_y[10367:10362] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1728 < i_size && h_count >= i_worm_x[10373:10368] * PIXEL_SIZE && h_count < i_worm_x[10373:10368] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10373:10368] * PIXEL_SIZE && v_count < i_worm_y[10373:10368] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1729 < i_size && h_count >= i_worm_x[10379:10374] * PIXEL_SIZE && h_count < i_worm_x[10379:10374] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10379:10374] * PIXEL_SIZE && v_count < i_worm_y[10379:10374] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1730 < i_size && h_count >= i_worm_x[10385:10380] * PIXEL_SIZE && h_count < i_worm_x[10385:10380] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10385:10380] * PIXEL_SIZE && v_count < i_worm_y[10385:10380] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1731 < i_size && h_count >= i_worm_x[10391:10386] * PIXEL_SIZE && h_count < i_worm_x[10391:10386] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10391:10386] * PIXEL_SIZE && v_count < i_worm_y[10391:10386] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1732 < i_size && h_count >= i_worm_x[10397:10392] * PIXEL_SIZE && h_count < i_worm_x[10397:10392] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10397:10392] * PIXEL_SIZE && v_count < i_worm_y[10397:10392] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1733 < i_size && h_count >= i_worm_x[10403:10398] * PIXEL_SIZE && h_count < i_worm_x[10403:10398] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10403:10398] * PIXEL_SIZE && v_count < i_worm_y[10403:10398] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1734 < i_size && h_count >= i_worm_x[10409:10404] * PIXEL_SIZE && h_count < i_worm_x[10409:10404] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10409:10404] * PIXEL_SIZE && v_count < i_worm_y[10409:10404] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1735 < i_size && h_count >= i_worm_x[10415:10410] * PIXEL_SIZE && h_count < i_worm_x[10415:10410] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10415:10410] * PIXEL_SIZE && v_count < i_worm_y[10415:10410] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1736 < i_size && h_count >= i_worm_x[10421:10416] * PIXEL_SIZE && h_count < i_worm_x[10421:10416] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10421:10416] * PIXEL_SIZE && v_count < i_worm_y[10421:10416] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1737 < i_size && h_count >= i_worm_x[10427:10422] * PIXEL_SIZE && h_count < i_worm_x[10427:10422] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10427:10422] * PIXEL_SIZE && v_count < i_worm_y[10427:10422] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1738 < i_size && h_count >= i_worm_x[10433:10428] * PIXEL_SIZE && h_count < i_worm_x[10433:10428] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10433:10428] * PIXEL_SIZE && v_count < i_worm_y[10433:10428] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1739 < i_size && h_count >= i_worm_x[10439:10434] * PIXEL_SIZE && h_count < i_worm_x[10439:10434] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10439:10434] * PIXEL_SIZE && v_count < i_worm_y[10439:10434] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1740 < i_size && h_count >= i_worm_x[10445:10440] * PIXEL_SIZE && h_count < i_worm_x[10445:10440] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10445:10440] * PIXEL_SIZE && v_count < i_worm_y[10445:10440] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1741 < i_size && h_count >= i_worm_x[10451:10446] * PIXEL_SIZE && h_count < i_worm_x[10451:10446] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10451:10446] * PIXEL_SIZE && v_count < i_worm_y[10451:10446] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1742 < i_size && h_count >= i_worm_x[10457:10452] * PIXEL_SIZE && h_count < i_worm_x[10457:10452] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10457:10452] * PIXEL_SIZE && v_count < i_worm_y[10457:10452] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1743 < i_size && h_count >= i_worm_x[10463:10458] * PIXEL_SIZE && h_count < i_worm_x[10463:10458] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10463:10458] * PIXEL_SIZE && v_count < i_worm_y[10463:10458] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1744 < i_size && h_count >= i_worm_x[10469:10464] * PIXEL_SIZE && h_count < i_worm_x[10469:10464] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10469:10464] * PIXEL_SIZE && v_count < i_worm_y[10469:10464] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1745 < i_size && h_count >= i_worm_x[10475:10470] * PIXEL_SIZE && h_count < i_worm_x[10475:10470] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10475:10470] * PIXEL_SIZE && v_count < i_worm_y[10475:10470] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1746 < i_size && h_count >= i_worm_x[10481:10476] * PIXEL_SIZE && h_count < i_worm_x[10481:10476] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10481:10476] * PIXEL_SIZE && v_count < i_worm_y[10481:10476] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1747 < i_size && h_count >= i_worm_x[10487:10482] * PIXEL_SIZE && h_count < i_worm_x[10487:10482] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10487:10482] * PIXEL_SIZE && v_count < i_worm_y[10487:10482] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1748 < i_size && h_count >= i_worm_x[10493:10488] * PIXEL_SIZE && h_count < i_worm_x[10493:10488] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10493:10488] * PIXEL_SIZE && v_count < i_worm_y[10493:10488] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1749 < i_size && h_count >= i_worm_x[10499:10494] * PIXEL_SIZE && h_count < i_worm_x[10499:10494] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10499:10494] * PIXEL_SIZE && v_count < i_worm_y[10499:10494] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1750 < i_size && h_count >= i_worm_x[10505:10500] * PIXEL_SIZE && h_count < i_worm_x[10505:10500] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10505:10500] * PIXEL_SIZE && v_count < i_worm_y[10505:10500] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1751 < i_size && h_count >= i_worm_x[10511:10506] * PIXEL_SIZE && h_count < i_worm_x[10511:10506] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10511:10506] * PIXEL_SIZE && v_count < i_worm_y[10511:10506] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1752 < i_size && h_count >= i_worm_x[10517:10512] * PIXEL_SIZE && h_count < i_worm_x[10517:10512] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10517:10512] * PIXEL_SIZE && v_count < i_worm_y[10517:10512] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1753 < i_size && h_count >= i_worm_x[10523:10518] * PIXEL_SIZE && h_count < i_worm_x[10523:10518] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10523:10518] * PIXEL_SIZE && v_count < i_worm_y[10523:10518] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1754 < i_size && h_count >= i_worm_x[10529:10524] * PIXEL_SIZE && h_count < i_worm_x[10529:10524] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10529:10524] * PIXEL_SIZE && v_count < i_worm_y[10529:10524] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1755 < i_size && h_count >= i_worm_x[10535:10530] * PIXEL_SIZE && h_count < i_worm_x[10535:10530] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10535:10530] * PIXEL_SIZE && v_count < i_worm_y[10535:10530] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1756 < i_size && h_count >= i_worm_x[10541:10536] * PIXEL_SIZE && h_count < i_worm_x[10541:10536] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10541:10536] * PIXEL_SIZE && v_count < i_worm_y[10541:10536] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1757 < i_size && h_count >= i_worm_x[10547:10542] * PIXEL_SIZE && h_count < i_worm_x[10547:10542] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10547:10542] * PIXEL_SIZE && v_count < i_worm_y[10547:10542] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1758 < i_size && h_count >= i_worm_x[10553:10548] * PIXEL_SIZE && h_count < i_worm_x[10553:10548] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10553:10548] * PIXEL_SIZE && v_count < i_worm_y[10553:10548] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1759 < i_size && h_count >= i_worm_x[10559:10554] * PIXEL_SIZE && h_count < i_worm_x[10559:10554] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10559:10554] * PIXEL_SIZE && v_count < i_worm_y[10559:10554] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1760 < i_size && h_count >= i_worm_x[10565:10560] * PIXEL_SIZE && h_count < i_worm_x[10565:10560] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10565:10560] * PIXEL_SIZE && v_count < i_worm_y[10565:10560] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1761 < i_size && h_count >= i_worm_x[10571:10566] * PIXEL_SIZE && h_count < i_worm_x[10571:10566] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10571:10566] * PIXEL_SIZE && v_count < i_worm_y[10571:10566] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1762 < i_size && h_count >= i_worm_x[10577:10572] * PIXEL_SIZE && h_count < i_worm_x[10577:10572] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10577:10572] * PIXEL_SIZE && v_count < i_worm_y[10577:10572] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1763 < i_size && h_count >= i_worm_x[10583:10578] * PIXEL_SIZE && h_count < i_worm_x[10583:10578] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10583:10578] * PIXEL_SIZE && v_count < i_worm_y[10583:10578] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1764 < i_size && h_count >= i_worm_x[10589:10584] * PIXEL_SIZE && h_count < i_worm_x[10589:10584] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10589:10584] * PIXEL_SIZE && v_count < i_worm_y[10589:10584] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1765 < i_size && h_count >= i_worm_x[10595:10590] * PIXEL_SIZE && h_count < i_worm_x[10595:10590] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10595:10590] * PIXEL_SIZE && v_count < i_worm_y[10595:10590] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1766 < i_size && h_count >= i_worm_x[10601:10596] * PIXEL_SIZE && h_count < i_worm_x[10601:10596] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10601:10596] * PIXEL_SIZE && v_count < i_worm_y[10601:10596] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1767 < i_size && h_count >= i_worm_x[10607:10602] * PIXEL_SIZE && h_count < i_worm_x[10607:10602] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10607:10602] * PIXEL_SIZE && v_count < i_worm_y[10607:10602] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1768 < i_size && h_count >= i_worm_x[10613:10608] * PIXEL_SIZE && h_count < i_worm_x[10613:10608] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10613:10608] * PIXEL_SIZE && v_count < i_worm_y[10613:10608] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1769 < i_size && h_count >= i_worm_x[10619:10614] * PIXEL_SIZE && h_count < i_worm_x[10619:10614] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10619:10614] * PIXEL_SIZE && v_count < i_worm_y[10619:10614] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1770 < i_size && h_count >= i_worm_x[10625:10620] * PIXEL_SIZE && h_count < i_worm_x[10625:10620] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10625:10620] * PIXEL_SIZE && v_count < i_worm_y[10625:10620] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1771 < i_size && h_count >= i_worm_x[10631:10626] * PIXEL_SIZE && h_count < i_worm_x[10631:10626] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10631:10626] * PIXEL_SIZE && v_count < i_worm_y[10631:10626] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1772 < i_size && h_count >= i_worm_x[10637:10632] * PIXEL_SIZE && h_count < i_worm_x[10637:10632] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10637:10632] * PIXEL_SIZE && v_count < i_worm_y[10637:10632] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1773 < i_size && h_count >= i_worm_x[10643:10638] * PIXEL_SIZE && h_count < i_worm_x[10643:10638] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10643:10638] * PIXEL_SIZE && v_count < i_worm_y[10643:10638] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1774 < i_size && h_count >= i_worm_x[10649:10644] * PIXEL_SIZE && h_count < i_worm_x[10649:10644] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10649:10644] * PIXEL_SIZE && v_count < i_worm_y[10649:10644] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1775 < i_size && h_count >= i_worm_x[10655:10650] * PIXEL_SIZE && h_count < i_worm_x[10655:10650] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10655:10650] * PIXEL_SIZE && v_count < i_worm_y[10655:10650] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1776 < i_size && h_count >= i_worm_x[10661:10656] * PIXEL_SIZE && h_count < i_worm_x[10661:10656] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10661:10656] * PIXEL_SIZE && v_count < i_worm_y[10661:10656] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1777 < i_size && h_count >= i_worm_x[10667:10662] * PIXEL_SIZE && h_count < i_worm_x[10667:10662] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10667:10662] * PIXEL_SIZE && v_count < i_worm_y[10667:10662] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1778 < i_size && h_count >= i_worm_x[10673:10668] * PIXEL_SIZE && h_count < i_worm_x[10673:10668] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10673:10668] * PIXEL_SIZE && v_count < i_worm_y[10673:10668] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1779 < i_size && h_count >= i_worm_x[10679:10674] * PIXEL_SIZE && h_count < i_worm_x[10679:10674] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10679:10674] * PIXEL_SIZE && v_count < i_worm_y[10679:10674] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1780 < i_size && h_count >= i_worm_x[10685:10680] * PIXEL_SIZE && h_count < i_worm_x[10685:10680] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10685:10680] * PIXEL_SIZE && v_count < i_worm_y[10685:10680] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1781 < i_size && h_count >= i_worm_x[10691:10686] * PIXEL_SIZE && h_count < i_worm_x[10691:10686] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10691:10686] * PIXEL_SIZE && v_count < i_worm_y[10691:10686] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1782 < i_size && h_count >= i_worm_x[10697:10692] * PIXEL_SIZE && h_count < i_worm_x[10697:10692] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10697:10692] * PIXEL_SIZE && v_count < i_worm_y[10697:10692] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1783 < i_size && h_count >= i_worm_x[10703:10698] * PIXEL_SIZE && h_count < i_worm_x[10703:10698] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10703:10698] * PIXEL_SIZE && v_count < i_worm_y[10703:10698] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1784 < i_size && h_count >= i_worm_x[10709:10704] * PIXEL_SIZE && h_count < i_worm_x[10709:10704] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10709:10704] * PIXEL_SIZE && v_count < i_worm_y[10709:10704] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1785 < i_size && h_count >= i_worm_x[10715:10710] * PIXEL_SIZE && h_count < i_worm_x[10715:10710] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10715:10710] * PIXEL_SIZE && v_count < i_worm_y[10715:10710] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1786 < i_size && h_count >= i_worm_x[10721:10716] * PIXEL_SIZE && h_count < i_worm_x[10721:10716] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10721:10716] * PIXEL_SIZE && v_count < i_worm_y[10721:10716] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1787 < i_size && h_count >= i_worm_x[10727:10722] * PIXEL_SIZE && h_count < i_worm_x[10727:10722] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10727:10722] * PIXEL_SIZE && v_count < i_worm_y[10727:10722] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1788 < i_size && h_count >= i_worm_x[10733:10728] * PIXEL_SIZE && h_count < i_worm_x[10733:10728] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10733:10728] * PIXEL_SIZE && v_count < i_worm_y[10733:10728] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1789 < i_size && h_count >= i_worm_x[10739:10734] * PIXEL_SIZE && h_count < i_worm_x[10739:10734] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10739:10734] * PIXEL_SIZE && v_count < i_worm_y[10739:10734] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1790 < i_size && h_count >= i_worm_x[10745:10740] * PIXEL_SIZE && h_count < i_worm_x[10745:10740] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10745:10740] * PIXEL_SIZE && v_count < i_worm_y[10745:10740] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1791 < i_size && h_count >= i_worm_x[10751:10746] * PIXEL_SIZE && h_count < i_worm_x[10751:10746] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10751:10746] * PIXEL_SIZE && v_count < i_worm_y[10751:10746] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1792 < i_size && h_count >= i_worm_x[10757:10752] * PIXEL_SIZE && h_count < i_worm_x[10757:10752] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10757:10752] * PIXEL_SIZE && v_count < i_worm_y[10757:10752] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1793 < i_size && h_count >= i_worm_x[10763:10758] * PIXEL_SIZE && h_count < i_worm_x[10763:10758] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10763:10758] * PIXEL_SIZE && v_count < i_worm_y[10763:10758] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1794 < i_size && h_count >= i_worm_x[10769:10764] * PIXEL_SIZE && h_count < i_worm_x[10769:10764] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10769:10764] * PIXEL_SIZE && v_count < i_worm_y[10769:10764] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1795 < i_size && h_count >= i_worm_x[10775:10770] * PIXEL_SIZE && h_count < i_worm_x[10775:10770] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10775:10770] * PIXEL_SIZE && v_count < i_worm_y[10775:10770] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1796 < i_size && h_count >= i_worm_x[10781:10776] * PIXEL_SIZE && h_count < i_worm_x[10781:10776] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10781:10776] * PIXEL_SIZE && v_count < i_worm_y[10781:10776] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1797 < i_size && h_count >= i_worm_x[10787:10782] * PIXEL_SIZE && h_count < i_worm_x[10787:10782] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10787:10782] * PIXEL_SIZE && v_count < i_worm_y[10787:10782] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1798 < i_size && h_count >= i_worm_x[10793:10788] * PIXEL_SIZE && h_count < i_worm_x[10793:10788] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10793:10788] * PIXEL_SIZE && v_count < i_worm_y[10793:10788] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1799 < i_size && h_count >= i_worm_x[10799:10794] * PIXEL_SIZE && h_count < i_worm_x[10799:10794] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10799:10794] * PIXEL_SIZE && v_count < i_worm_y[10799:10794] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1800 < i_size && h_count >= i_worm_x[10805:10800] * PIXEL_SIZE && h_count < i_worm_x[10805:10800] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10805:10800] * PIXEL_SIZE && v_count < i_worm_y[10805:10800] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1801 < i_size && h_count >= i_worm_x[10811:10806] * PIXEL_SIZE && h_count < i_worm_x[10811:10806] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10811:10806] * PIXEL_SIZE && v_count < i_worm_y[10811:10806] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1802 < i_size && h_count >= i_worm_x[10817:10812] * PIXEL_SIZE && h_count < i_worm_x[10817:10812] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10817:10812] * PIXEL_SIZE && v_count < i_worm_y[10817:10812] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1803 < i_size && h_count >= i_worm_x[10823:10818] * PIXEL_SIZE && h_count < i_worm_x[10823:10818] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10823:10818] * PIXEL_SIZE && v_count < i_worm_y[10823:10818] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1804 < i_size && h_count >= i_worm_x[10829:10824] * PIXEL_SIZE && h_count < i_worm_x[10829:10824] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10829:10824] * PIXEL_SIZE && v_count < i_worm_y[10829:10824] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1805 < i_size && h_count >= i_worm_x[10835:10830] * PIXEL_SIZE && h_count < i_worm_x[10835:10830] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10835:10830] * PIXEL_SIZE && v_count < i_worm_y[10835:10830] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1806 < i_size && h_count >= i_worm_x[10841:10836] * PIXEL_SIZE && h_count < i_worm_x[10841:10836] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10841:10836] * PIXEL_SIZE && v_count < i_worm_y[10841:10836] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1807 < i_size && h_count >= i_worm_x[10847:10842] * PIXEL_SIZE && h_count < i_worm_x[10847:10842] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10847:10842] * PIXEL_SIZE && v_count < i_worm_y[10847:10842] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1808 < i_size && h_count >= i_worm_x[10853:10848] * PIXEL_SIZE && h_count < i_worm_x[10853:10848] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10853:10848] * PIXEL_SIZE && v_count < i_worm_y[10853:10848] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1809 < i_size && h_count >= i_worm_x[10859:10854] * PIXEL_SIZE && h_count < i_worm_x[10859:10854] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10859:10854] * PIXEL_SIZE && v_count < i_worm_y[10859:10854] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1810 < i_size && h_count >= i_worm_x[10865:10860] * PIXEL_SIZE && h_count < i_worm_x[10865:10860] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10865:10860] * PIXEL_SIZE && v_count < i_worm_y[10865:10860] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1811 < i_size && h_count >= i_worm_x[10871:10866] * PIXEL_SIZE && h_count < i_worm_x[10871:10866] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10871:10866] * PIXEL_SIZE && v_count < i_worm_y[10871:10866] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1812 < i_size && h_count >= i_worm_x[10877:10872] * PIXEL_SIZE && h_count < i_worm_x[10877:10872] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10877:10872] * PIXEL_SIZE && v_count < i_worm_y[10877:10872] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1813 < i_size && h_count >= i_worm_x[10883:10878] * PIXEL_SIZE && h_count < i_worm_x[10883:10878] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10883:10878] * PIXEL_SIZE && v_count < i_worm_y[10883:10878] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1814 < i_size && h_count >= i_worm_x[10889:10884] * PIXEL_SIZE && h_count < i_worm_x[10889:10884] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10889:10884] * PIXEL_SIZE && v_count < i_worm_y[10889:10884] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1815 < i_size && h_count >= i_worm_x[10895:10890] * PIXEL_SIZE && h_count < i_worm_x[10895:10890] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10895:10890] * PIXEL_SIZE && v_count < i_worm_y[10895:10890] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1816 < i_size && h_count >= i_worm_x[10901:10896] * PIXEL_SIZE && h_count < i_worm_x[10901:10896] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10901:10896] * PIXEL_SIZE && v_count < i_worm_y[10901:10896] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1817 < i_size && h_count >= i_worm_x[10907:10902] * PIXEL_SIZE && h_count < i_worm_x[10907:10902] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10907:10902] * PIXEL_SIZE && v_count < i_worm_y[10907:10902] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1818 < i_size && h_count >= i_worm_x[10913:10908] * PIXEL_SIZE && h_count < i_worm_x[10913:10908] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10913:10908] * PIXEL_SIZE && v_count < i_worm_y[10913:10908] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1819 < i_size && h_count >= i_worm_x[10919:10914] * PIXEL_SIZE && h_count < i_worm_x[10919:10914] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10919:10914] * PIXEL_SIZE && v_count < i_worm_y[10919:10914] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1820 < i_size && h_count >= i_worm_x[10925:10920] * PIXEL_SIZE && h_count < i_worm_x[10925:10920] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10925:10920] * PIXEL_SIZE && v_count < i_worm_y[10925:10920] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1821 < i_size && h_count >= i_worm_x[10931:10926] * PIXEL_SIZE && h_count < i_worm_x[10931:10926] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10931:10926] * PIXEL_SIZE && v_count < i_worm_y[10931:10926] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1822 < i_size && h_count >= i_worm_x[10937:10932] * PIXEL_SIZE && h_count < i_worm_x[10937:10932] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10937:10932] * PIXEL_SIZE && v_count < i_worm_y[10937:10932] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1823 < i_size && h_count >= i_worm_x[10943:10938] * PIXEL_SIZE && h_count < i_worm_x[10943:10938] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10943:10938] * PIXEL_SIZE && v_count < i_worm_y[10943:10938] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1824 < i_size && h_count >= i_worm_x[10949:10944] * PIXEL_SIZE && h_count < i_worm_x[10949:10944] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10949:10944] * PIXEL_SIZE && v_count < i_worm_y[10949:10944] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1825 < i_size && h_count >= i_worm_x[10955:10950] * PIXEL_SIZE && h_count < i_worm_x[10955:10950] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10955:10950] * PIXEL_SIZE && v_count < i_worm_y[10955:10950] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1826 < i_size && h_count >= i_worm_x[10961:10956] * PIXEL_SIZE && h_count < i_worm_x[10961:10956] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10961:10956] * PIXEL_SIZE && v_count < i_worm_y[10961:10956] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1827 < i_size && h_count >= i_worm_x[10967:10962] * PIXEL_SIZE && h_count < i_worm_x[10967:10962] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10967:10962] * PIXEL_SIZE && v_count < i_worm_y[10967:10962] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1828 < i_size && h_count >= i_worm_x[10973:10968] * PIXEL_SIZE && h_count < i_worm_x[10973:10968] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10973:10968] * PIXEL_SIZE && v_count < i_worm_y[10973:10968] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1829 < i_size && h_count >= i_worm_x[10979:10974] * PIXEL_SIZE && h_count < i_worm_x[10979:10974] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10979:10974] * PIXEL_SIZE && v_count < i_worm_y[10979:10974] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1830 < i_size && h_count >= i_worm_x[10985:10980] * PIXEL_SIZE && h_count < i_worm_x[10985:10980] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10985:10980] * PIXEL_SIZE && v_count < i_worm_y[10985:10980] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1831 < i_size && h_count >= i_worm_x[10991:10986] * PIXEL_SIZE && h_count < i_worm_x[10991:10986] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10991:10986] * PIXEL_SIZE && v_count < i_worm_y[10991:10986] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1832 < i_size && h_count >= i_worm_x[10997:10992] * PIXEL_SIZE && h_count < i_worm_x[10997:10992] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[10997:10992] * PIXEL_SIZE && v_count < i_worm_y[10997:10992] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1833 < i_size && h_count >= i_worm_x[11003:10998] * PIXEL_SIZE && h_count < i_worm_x[11003:10998] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11003:10998] * PIXEL_SIZE && v_count < i_worm_y[11003:10998] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1834 < i_size && h_count >= i_worm_x[11009:11004] * PIXEL_SIZE && h_count < i_worm_x[11009:11004] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11009:11004] * PIXEL_SIZE && v_count < i_worm_y[11009:11004] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1835 < i_size && h_count >= i_worm_x[11015:11010] * PIXEL_SIZE && h_count < i_worm_x[11015:11010] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11015:11010] * PIXEL_SIZE && v_count < i_worm_y[11015:11010] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1836 < i_size && h_count >= i_worm_x[11021:11016] * PIXEL_SIZE && h_count < i_worm_x[11021:11016] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11021:11016] * PIXEL_SIZE && v_count < i_worm_y[11021:11016] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1837 < i_size && h_count >= i_worm_x[11027:11022] * PIXEL_SIZE && h_count < i_worm_x[11027:11022] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11027:11022] * PIXEL_SIZE && v_count < i_worm_y[11027:11022] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1838 < i_size && h_count >= i_worm_x[11033:11028] * PIXEL_SIZE && h_count < i_worm_x[11033:11028] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11033:11028] * PIXEL_SIZE && v_count < i_worm_y[11033:11028] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1839 < i_size && h_count >= i_worm_x[11039:11034] * PIXEL_SIZE && h_count < i_worm_x[11039:11034] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11039:11034] * PIXEL_SIZE && v_count < i_worm_y[11039:11034] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1840 < i_size && h_count >= i_worm_x[11045:11040] * PIXEL_SIZE && h_count < i_worm_x[11045:11040] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11045:11040] * PIXEL_SIZE && v_count < i_worm_y[11045:11040] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1841 < i_size && h_count >= i_worm_x[11051:11046] * PIXEL_SIZE && h_count < i_worm_x[11051:11046] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11051:11046] * PIXEL_SIZE && v_count < i_worm_y[11051:11046] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1842 < i_size && h_count >= i_worm_x[11057:11052] * PIXEL_SIZE && h_count < i_worm_x[11057:11052] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11057:11052] * PIXEL_SIZE && v_count < i_worm_y[11057:11052] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1843 < i_size && h_count >= i_worm_x[11063:11058] * PIXEL_SIZE && h_count < i_worm_x[11063:11058] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11063:11058] * PIXEL_SIZE && v_count < i_worm_y[11063:11058] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1844 < i_size && h_count >= i_worm_x[11069:11064] * PIXEL_SIZE && h_count < i_worm_x[11069:11064] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11069:11064] * PIXEL_SIZE && v_count < i_worm_y[11069:11064] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1845 < i_size && h_count >= i_worm_x[11075:11070] * PIXEL_SIZE && h_count < i_worm_x[11075:11070] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11075:11070] * PIXEL_SIZE && v_count < i_worm_y[11075:11070] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1846 < i_size && h_count >= i_worm_x[11081:11076] * PIXEL_SIZE && h_count < i_worm_x[11081:11076] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11081:11076] * PIXEL_SIZE && v_count < i_worm_y[11081:11076] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1847 < i_size && h_count >= i_worm_x[11087:11082] * PIXEL_SIZE && h_count < i_worm_x[11087:11082] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11087:11082] * PIXEL_SIZE && v_count < i_worm_y[11087:11082] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1848 < i_size && h_count >= i_worm_x[11093:11088] * PIXEL_SIZE && h_count < i_worm_x[11093:11088] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11093:11088] * PIXEL_SIZE && v_count < i_worm_y[11093:11088] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1849 < i_size && h_count >= i_worm_x[11099:11094] * PIXEL_SIZE && h_count < i_worm_x[11099:11094] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11099:11094] * PIXEL_SIZE && v_count < i_worm_y[11099:11094] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1850 < i_size && h_count >= i_worm_x[11105:11100] * PIXEL_SIZE && h_count < i_worm_x[11105:11100] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11105:11100] * PIXEL_SIZE && v_count < i_worm_y[11105:11100] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1851 < i_size && h_count >= i_worm_x[11111:11106] * PIXEL_SIZE && h_count < i_worm_x[11111:11106] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11111:11106] * PIXEL_SIZE && v_count < i_worm_y[11111:11106] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1852 < i_size && h_count >= i_worm_x[11117:11112] * PIXEL_SIZE && h_count < i_worm_x[11117:11112] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11117:11112] * PIXEL_SIZE && v_count < i_worm_y[11117:11112] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1853 < i_size && h_count >= i_worm_x[11123:11118] * PIXEL_SIZE && h_count < i_worm_x[11123:11118] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11123:11118] * PIXEL_SIZE && v_count < i_worm_y[11123:11118] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1854 < i_size && h_count >= i_worm_x[11129:11124] * PIXEL_SIZE && h_count < i_worm_x[11129:11124] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11129:11124] * PIXEL_SIZE && v_count < i_worm_y[11129:11124] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1855 < i_size && h_count >= i_worm_x[11135:11130] * PIXEL_SIZE && h_count < i_worm_x[11135:11130] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11135:11130] * PIXEL_SIZE && v_count < i_worm_y[11135:11130] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1856 < i_size && h_count >= i_worm_x[11141:11136] * PIXEL_SIZE && h_count < i_worm_x[11141:11136] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11141:11136] * PIXEL_SIZE && v_count < i_worm_y[11141:11136] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1857 < i_size && h_count >= i_worm_x[11147:11142] * PIXEL_SIZE && h_count < i_worm_x[11147:11142] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11147:11142] * PIXEL_SIZE && v_count < i_worm_y[11147:11142] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1858 < i_size && h_count >= i_worm_x[11153:11148] * PIXEL_SIZE && h_count < i_worm_x[11153:11148] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11153:11148] * PIXEL_SIZE && v_count < i_worm_y[11153:11148] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1859 < i_size && h_count >= i_worm_x[11159:11154] * PIXEL_SIZE && h_count < i_worm_x[11159:11154] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11159:11154] * PIXEL_SIZE && v_count < i_worm_y[11159:11154] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1860 < i_size && h_count >= i_worm_x[11165:11160] * PIXEL_SIZE && h_count < i_worm_x[11165:11160] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11165:11160] * PIXEL_SIZE && v_count < i_worm_y[11165:11160] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1861 < i_size && h_count >= i_worm_x[11171:11166] * PIXEL_SIZE && h_count < i_worm_x[11171:11166] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11171:11166] * PIXEL_SIZE && v_count < i_worm_y[11171:11166] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1862 < i_size && h_count >= i_worm_x[11177:11172] * PIXEL_SIZE && h_count < i_worm_x[11177:11172] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11177:11172] * PIXEL_SIZE && v_count < i_worm_y[11177:11172] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1863 < i_size && h_count >= i_worm_x[11183:11178] * PIXEL_SIZE && h_count < i_worm_x[11183:11178] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11183:11178] * PIXEL_SIZE && v_count < i_worm_y[11183:11178] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1864 < i_size && h_count >= i_worm_x[11189:11184] * PIXEL_SIZE && h_count < i_worm_x[11189:11184] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11189:11184] * PIXEL_SIZE && v_count < i_worm_y[11189:11184] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1865 < i_size && h_count >= i_worm_x[11195:11190] * PIXEL_SIZE && h_count < i_worm_x[11195:11190] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11195:11190] * PIXEL_SIZE && v_count < i_worm_y[11195:11190] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1866 < i_size && h_count >= i_worm_x[11201:11196] * PIXEL_SIZE && h_count < i_worm_x[11201:11196] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11201:11196] * PIXEL_SIZE && v_count < i_worm_y[11201:11196] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1867 < i_size && h_count >= i_worm_x[11207:11202] * PIXEL_SIZE && h_count < i_worm_x[11207:11202] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11207:11202] * PIXEL_SIZE && v_count < i_worm_y[11207:11202] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1868 < i_size && h_count >= i_worm_x[11213:11208] * PIXEL_SIZE && h_count < i_worm_x[11213:11208] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11213:11208] * PIXEL_SIZE && v_count < i_worm_y[11213:11208] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1869 < i_size && h_count >= i_worm_x[11219:11214] * PIXEL_SIZE && h_count < i_worm_x[11219:11214] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11219:11214] * PIXEL_SIZE && v_count < i_worm_y[11219:11214] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1870 < i_size && h_count >= i_worm_x[11225:11220] * PIXEL_SIZE && h_count < i_worm_x[11225:11220] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11225:11220] * PIXEL_SIZE && v_count < i_worm_y[11225:11220] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1871 < i_size && h_count >= i_worm_x[11231:11226] * PIXEL_SIZE && h_count < i_worm_x[11231:11226] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11231:11226] * PIXEL_SIZE && v_count < i_worm_y[11231:11226] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1872 < i_size && h_count >= i_worm_x[11237:11232] * PIXEL_SIZE && h_count < i_worm_x[11237:11232] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11237:11232] * PIXEL_SIZE && v_count < i_worm_y[11237:11232] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1873 < i_size && h_count >= i_worm_x[11243:11238] * PIXEL_SIZE && h_count < i_worm_x[11243:11238] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11243:11238] * PIXEL_SIZE && v_count < i_worm_y[11243:11238] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1874 < i_size && h_count >= i_worm_x[11249:11244] * PIXEL_SIZE && h_count < i_worm_x[11249:11244] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11249:11244] * PIXEL_SIZE && v_count < i_worm_y[11249:11244] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1875 < i_size && h_count >= i_worm_x[11255:11250] * PIXEL_SIZE && h_count < i_worm_x[11255:11250] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11255:11250] * PIXEL_SIZE && v_count < i_worm_y[11255:11250] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1876 < i_size && h_count >= i_worm_x[11261:11256] * PIXEL_SIZE && h_count < i_worm_x[11261:11256] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11261:11256] * PIXEL_SIZE && v_count < i_worm_y[11261:11256] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1877 < i_size && h_count >= i_worm_x[11267:11262] * PIXEL_SIZE && h_count < i_worm_x[11267:11262] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11267:11262] * PIXEL_SIZE && v_count < i_worm_y[11267:11262] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1878 < i_size && h_count >= i_worm_x[11273:11268] * PIXEL_SIZE && h_count < i_worm_x[11273:11268] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11273:11268] * PIXEL_SIZE && v_count < i_worm_y[11273:11268] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1879 < i_size && h_count >= i_worm_x[11279:11274] * PIXEL_SIZE && h_count < i_worm_x[11279:11274] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11279:11274] * PIXEL_SIZE && v_count < i_worm_y[11279:11274] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1880 < i_size && h_count >= i_worm_x[11285:11280] * PIXEL_SIZE && h_count < i_worm_x[11285:11280] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11285:11280] * PIXEL_SIZE && v_count < i_worm_y[11285:11280] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1881 < i_size && h_count >= i_worm_x[11291:11286] * PIXEL_SIZE && h_count < i_worm_x[11291:11286] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11291:11286] * PIXEL_SIZE && v_count < i_worm_y[11291:11286] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1882 < i_size && h_count >= i_worm_x[11297:11292] * PIXEL_SIZE && h_count < i_worm_x[11297:11292] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11297:11292] * PIXEL_SIZE && v_count < i_worm_y[11297:11292] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1883 < i_size && h_count >= i_worm_x[11303:11298] * PIXEL_SIZE && h_count < i_worm_x[11303:11298] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11303:11298] * PIXEL_SIZE && v_count < i_worm_y[11303:11298] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1884 < i_size && h_count >= i_worm_x[11309:11304] * PIXEL_SIZE && h_count < i_worm_x[11309:11304] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11309:11304] * PIXEL_SIZE && v_count < i_worm_y[11309:11304] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1885 < i_size && h_count >= i_worm_x[11315:11310] * PIXEL_SIZE && h_count < i_worm_x[11315:11310] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11315:11310] * PIXEL_SIZE && v_count < i_worm_y[11315:11310] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1886 < i_size && h_count >= i_worm_x[11321:11316] * PIXEL_SIZE && h_count < i_worm_x[11321:11316] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11321:11316] * PIXEL_SIZE && v_count < i_worm_y[11321:11316] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1887 < i_size && h_count >= i_worm_x[11327:11322] * PIXEL_SIZE && h_count < i_worm_x[11327:11322] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11327:11322] * PIXEL_SIZE && v_count < i_worm_y[11327:11322] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1888 < i_size && h_count >= i_worm_x[11333:11328] * PIXEL_SIZE && h_count < i_worm_x[11333:11328] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11333:11328] * PIXEL_SIZE && v_count < i_worm_y[11333:11328] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1889 < i_size && h_count >= i_worm_x[11339:11334] * PIXEL_SIZE && h_count < i_worm_x[11339:11334] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11339:11334] * PIXEL_SIZE && v_count < i_worm_y[11339:11334] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1890 < i_size && h_count >= i_worm_x[11345:11340] * PIXEL_SIZE && h_count < i_worm_x[11345:11340] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11345:11340] * PIXEL_SIZE && v_count < i_worm_y[11345:11340] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1891 < i_size && h_count >= i_worm_x[11351:11346] * PIXEL_SIZE && h_count < i_worm_x[11351:11346] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11351:11346] * PIXEL_SIZE && v_count < i_worm_y[11351:11346] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1892 < i_size && h_count >= i_worm_x[11357:11352] * PIXEL_SIZE && h_count < i_worm_x[11357:11352] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11357:11352] * PIXEL_SIZE && v_count < i_worm_y[11357:11352] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1893 < i_size && h_count >= i_worm_x[11363:11358] * PIXEL_SIZE && h_count < i_worm_x[11363:11358] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11363:11358] * PIXEL_SIZE && v_count < i_worm_y[11363:11358] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1894 < i_size && h_count >= i_worm_x[11369:11364] * PIXEL_SIZE && h_count < i_worm_x[11369:11364] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11369:11364] * PIXEL_SIZE && v_count < i_worm_y[11369:11364] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1895 < i_size && h_count >= i_worm_x[11375:11370] * PIXEL_SIZE && h_count < i_worm_x[11375:11370] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11375:11370] * PIXEL_SIZE && v_count < i_worm_y[11375:11370] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1896 < i_size && h_count >= i_worm_x[11381:11376] * PIXEL_SIZE && h_count < i_worm_x[11381:11376] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11381:11376] * PIXEL_SIZE && v_count < i_worm_y[11381:11376] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1897 < i_size && h_count >= i_worm_x[11387:11382] * PIXEL_SIZE && h_count < i_worm_x[11387:11382] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11387:11382] * PIXEL_SIZE && v_count < i_worm_y[11387:11382] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1898 < i_size && h_count >= i_worm_x[11393:11388] * PIXEL_SIZE && h_count < i_worm_x[11393:11388] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11393:11388] * PIXEL_SIZE && v_count < i_worm_y[11393:11388] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1899 < i_size && h_count >= i_worm_x[11399:11394] * PIXEL_SIZE && h_count < i_worm_x[11399:11394] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11399:11394] * PIXEL_SIZE && v_count < i_worm_y[11399:11394] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1900 < i_size && h_count >= i_worm_x[11405:11400] * PIXEL_SIZE && h_count < i_worm_x[11405:11400] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11405:11400] * PIXEL_SIZE && v_count < i_worm_y[11405:11400] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1901 < i_size && h_count >= i_worm_x[11411:11406] * PIXEL_SIZE && h_count < i_worm_x[11411:11406] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11411:11406] * PIXEL_SIZE && v_count < i_worm_y[11411:11406] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1902 < i_size && h_count >= i_worm_x[11417:11412] * PIXEL_SIZE && h_count < i_worm_x[11417:11412] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11417:11412] * PIXEL_SIZE && v_count < i_worm_y[11417:11412] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1903 < i_size && h_count >= i_worm_x[11423:11418] * PIXEL_SIZE && h_count < i_worm_x[11423:11418] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11423:11418] * PIXEL_SIZE && v_count < i_worm_y[11423:11418] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1904 < i_size && h_count >= i_worm_x[11429:11424] * PIXEL_SIZE && h_count < i_worm_x[11429:11424] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11429:11424] * PIXEL_SIZE && v_count < i_worm_y[11429:11424] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1905 < i_size && h_count >= i_worm_x[11435:11430] * PIXEL_SIZE && h_count < i_worm_x[11435:11430] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11435:11430] * PIXEL_SIZE && v_count < i_worm_y[11435:11430] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1906 < i_size && h_count >= i_worm_x[11441:11436] * PIXEL_SIZE && h_count < i_worm_x[11441:11436] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11441:11436] * PIXEL_SIZE && v_count < i_worm_y[11441:11436] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1907 < i_size && h_count >= i_worm_x[11447:11442] * PIXEL_SIZE && h_count < i_worm_x[11447:11442] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11447:11442] * PIXEL_SIZE && v_count < i_worm_y[11447:11442] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1908 < i_size && h_count >= i_worm_x[11453:11448] * PIXEL_SIZE && h_count < i_worm_x[11453:11448] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11453:11448] * PIXEL_SIZE && v_count < i_worm_y[11453:11448] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1909 < i_size && h_count >= i_worm_x[11459:11454] * PIXEL_SIZE && h_count < i_worm_x[11459:11454] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11459:11454] * PIXEL_SIZE && v_count < i_worm_y[11459:11454] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1910 < i_size && h_count >= i_worm_x[11465:11460] * PIXEL_SIZE && h_count < i_worm_x[11465:11460] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11465:11460] * PIXEL_SIZE && v_count < i_worm_y[11465:11460] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1911 < i_size && h_count >= i_worm_x[11471:11466] * PIXEL_SIZE && h_count < i_worm_x[11471:11466] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11471:11466] * PIXEL_SIZE && v_count < i_worm_y[11471:11466] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1912 < i_size && h_count >= i_worm_x[11477:11472] * PIXEL_SIZE && h_count < i_worm_x[11477:11472] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11477:11472] * PIXEL_SIZE && v_count < i_worm_y[11477:11472] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1913 < i_size && h_count >= i_worm_x[11483:11478] * PIXEL_SIZE && h_count < i_worm_x[11483:11478] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11483:11478] * PIXEL_SIZE && v_count < i_worm_y[11483:11478] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1914 < i_size && h_count >= i_worm_x[11489:11484] * PIXEL_SIZE && h_count < i_worm_x[11489:11484] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11489:11484] * PIXEL_SIZE && v_count < i_worm_y[11489:11484] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1915 < i_size && h_count >= i_worm_x[11495:11490] * PIXEL_SIZE && h_count < i_worm_x[11495:11490] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11495:11490] * PIXEL_SIZE && v_count < i_worm_y[11495:11490] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1916 < i_size && h_count >= i_worm_x[11501:11496] * PIXEL_SIZE && h_count < i_worm_x[11501:11496] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11501:11496] * PIXEL_SIZE && v_count < i_worm_y[11501:11496] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1917 < i_size && h_count >= i_worm_x[11507:11502] * PIXEL_SIZE && h_count < i_worm_x[11507:11502] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11507:11502] * PIXEL_SIZE && v_count < i_worm_y[11507:11502] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1918 < i_size && h_count >= i_worm_x[11513:11508] * PIXEL_SIZE && h_count < i_worm_x[11513:11508] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11513:11508] * PIXEL_SIZE && v_count < i_worm_y[11513:11508] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1919 < i_size && h_count >= i_worm_x[11519:11514] * PIXEL_SIZE && h_count < i_worm_x[11519:11514] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11519:11514] * PIXEL_SIZE && v_count < i_worm_y[11519:11514] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1920 < i_size && h_count >= i_worm_x[11525:11520] * PIXEL_SIZE && h_count < i_worm_x[11525:11520] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11525:11520] * PIXEL_SIZE && v_count < i_worm_y[11525:11520] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1921 < i_size && h_count >= i_worm_x[11531:11526] * PIXEL_SIZE && h_count < i_worm_x[11531:11526] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11531:11526] * PIXEL_SIZE && v_count < i_worm_y[11531:11526] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1922 < i_size && h_count >= i_worm_x[11537:11532] * PIXEL_SIZE && h_count < i_worm_x[11537:11532] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11537:11532] * PIXEL_SIZE && v_count < i_worm_y[11537:11532] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1923 < i_size && h_count >= i_worm_x[11543:11538] * PIXEL_SIZE && h_count < i_worm_x[11543:11538] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11543:11538] * PIXEL_SIZE && v_count < i_worm_y[11543:11538] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1924 < i_size && h_count >= i_worm_x[11549:11544] * PIXEL_SIZE && h_count < i_worm_x[11549:11544] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11549:11544] * PIXEL_SIZE && v_count < i_worm_y[11549:11544] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1925 < i_size && h_count >= i_worm_x[11555:11550] * PIXEL_SIZE && h_count < i_worm_x[11555:11550] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11555:11550] * PIXEL_SIZE && v_count < i_worm_y[11555:11550] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1926 < i_size && h_count >= i_worm_x[11561:11556] * PIXEL_SIZE && h_count < i_worm_x[11561:11556] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11561:11556] * PIXEL_SIZE && v_count < i_worm_y[11561:11556] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1927 < i_size && h_count >= i_worm_x[11567:11562] * PIXEL_SIZE && h_count < i_worm_x[11567:11562] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11567:11562] * PIXEL_SIZE && v_count < i_worm_y[11567:11562] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1928 < i_size && h_count >= i_worm_x[11573:11568] * PIXEL_SIZE && h_count < i_worm_x[11573:11568] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11573:11568] * PIXEL_SIZE && v_count < i_worm_y[11573:11568] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1929 < i_size && h_count >= i_worm_x[11579:11574] * PIXEL_SIZE && h_count < i_worm_x[11579:11574] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11579:11574] * PIXEL_SIZE && v_count < i_worm_y[11579:11574] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1930 < i_size && h_count >= i_worm_x[11585:11580] * PIXEL_SIZE && h_count < i_worm_x[11585:11580] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11585:11580] * PIXEL_SIZE && v_count < i_worm_y[11585:11580] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1931 < i_size && h_count >= i_worm_x[11591:11586] * PIXEL_SIZE && h_count < i_worm_x[11591:11586] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11591:11586] * PIXEL_SIZE && v_count < i_worm_y[11591:11586] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1932 < i_size && h_count >= i_worm_x[11597:11592] * PIXEL_SIZE && h_count < i_worm_x[11597:11592] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11597:11592] * PIXEL_SIZE && v_count < i_worm_y[11597:11592] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1933 < i_size && h_count >= i_worm_x[11603:11598] * PIXEL_SIZE && h_count < i_worm_x[11603:11598] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11603:11598] * PIXEL_SIZE && v_count < i_worm_y[11603:11598] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1934 < i_size && h_count >= i_worm_x[11609:11604] * PIXEL_SIZE && h_count < i_worm_x[11609:11604] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11609:11604] * PIXEL_SIZE && v_count < i_worm_y[11609:11604] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1935 < i_size && h_count >= i_worm_x[11615:11610] * PIXEL_SIZE && h_count < i_worm_x[11615:11610] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11615:11610] * PIXEL_SIZE && v_count < i_worm_y[11615:11610] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1936 < i_size && h_count >= i_worm_x[11621:11616] * PIXEL_SIZE && h_count < i_worm_x[11621:11616] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11621:11616] * PIXEL_SIZE && v_count < i_worm_y[11621:11616] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1937 < i_size && h_count >= i_worm_x[11627:11622] * PIXEL_SIZE && h_count < i_worm_x[11627:11622] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11627:11622] * PIXEL_SIZE && v_count < i_worm_y[11627:11622] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1938 < i_size && h_count >= i_worm_x[11633:11628] * PIXEL_SIZE && h_count < i_worm_x[11633:11628] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11633:11628] * PIXEL_SIZE && v_count < i_worm_y[11633:11628] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1939 < i_size && h_count >= i_worm_x[11639:11634] * PIXEL_SIZE && h_count < i_worm_x[11639:11634] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11639:11634] * PIXEL_SIZE && v_count < i_worm_y[11639:11634] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1940 < i_size && h_count >= i_worm_x[11645:11640] * PIXEL_SIZE && h_count < i_worm_x[11645:11640] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11645:11640] * PIXEL_SIZE && v_count < i_worm_y[11645:11640] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1941 < i_size && h_count >= i_worm_x[11651:11646] * PIXEL_SIZE && h_count < i_worm_x[11651:11646] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11651:11646] * PIXEL_SIZE && v_count < i_worm_y[11651:11646] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1942 < i_size && h_count >= i_worm_x[11657:11652] * PIXEL_SIZE && h_count < i_worm_x[11657:11652] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11657:11652] * PIXEL_SIZE && v_count < i_worm_y[11657:11652] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1943 < i_size && h_count >= i_worm_x[11663:11658] * PIXEL_SIZE && h_count < i_worm_x[11663:11658] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11663:11658] * PIXEL_SIZE && v_count < i_worm_y[11663:11658] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1944 < i_size && h_count >= i_worm_x[11669:11664] * PIXEL_SIZE && h_count < i_worm_x[11669:11664] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11669:11664] * PIXEL_SIZE && v_count < i_worm_y[11669:11664] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1945 < i_size && h_count >= i_worm_x[11675:11670] * PIXEL_SIZE && h_count < i_worm_x[11675:11670] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11675:11670] * PIXEL_SIZE && v_count < i_worm_y[11675:11670] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1946 < i_size && h_count >= i_worm_x[11681:11676] * PIXEL_SIZE && h_count < i_worm_x[11681:11676] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11681:11676] * PIXEL_SIZE && v_count < i_worm_y[11681:11676] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1947 < i_size && h_count >= i_worm_x[11687:11682] * PIXEL_SIZE && h_count < i_worm_x[11687:11682] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11687:11682] * PIXEL_SIZE && v_count < i_worm_y[11687:11682] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1948 < i_size && h_count >= i_worm_x[11693:11688] * PIXEL_SIZE && h_count < i_worm_x[11693:11688] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11693:11688] * PIXEL_SIZE && v_count < i_worm_y[11693:11688] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1949 < i_size && h_count >= i_worm_x[11699:11694] * PIXEL_SIZE && h_count < i_worm_x[11699:11694] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11699:11694] * PIXEL_SIZE && v_count < i_worm_y[11699:11694] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1950 < i_size && h_count >= i_worm_x[11705:11700] * PIXEL_SIZE && h_count < i_worm_x[11705:11700] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11705:11700] * PIXEL_SIZE && v_count < i_worm_y[11705:11700] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1951 < i_size && h_count >= i_worm_x[11711:11706] * PIXEL_SIZE && h_count < i_worm_x[11711:11706] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11711:11706] * PIXEL_SIZE && v_count < i_worm_y[11711:11706] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1952 < i_size && h_count >= i_worm_x[11717:11712] * PIXEL_SIZE && h_count < i_worm_x[11717:11712] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11717:11712] * PIXEL_SIZE && v_count < i_worm_y[11717:11712] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1953 < i_size && h_count >= i_worm_x[11723:11718] * PIXEL_SIZE && h_count < i_worm_x[11723:11718] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11723:11718] * PIXEL_SIZE && v_count < i_worm_y[11723:11718] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1954 < i_size && h_count >= i_worm_x[11729:11724] * PIXEL_SIZE && h_count < i_worm_x[11729:11724] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11729:11724] * PIXEL_SIZE && v_count < i_worm_y[11729:11724] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1955 < i_size && h_count >= i_worm_x[11735:11730] * PIXEL_SIZE && h_count < i_worm_x[11735:11730] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11735:11730] * PIXEL_SIZE && v_count < i_worm_y[11735:11730] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1956 < i_size && h_count >= i_worm_x[11741:11736] * PIXEL_SIZE && h_count < i_worm_x[11741:11736] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11741:11736] * PIXEL_SIZE && v_count < i_worm_y[11741:11736] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1957 < i_size && h_count >= i_worm_x[11747:11742] * PIXEL_SIZE && h_count < i_worm_x[11747:11742] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11747:11742] * PIXEL_SIZE && v_count < i_worm_y[11747:11742] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1958 < i_size && h_count >= i_worm_x[11753:11748] * PIXEL_SIZE && h_count < i_worm_x[11753:11748] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11753:11748] * PIXEL_SIZE && v_count < i_worm_y[11753:11748] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1959 < i_size && h_count >= i_worm_x[11759:11754] * PIXEL_SIZE && h_count < i_worm_x[11759:11754] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11759:11754] * PIXEL_SIZE && v_count < i_worm_y[11759:11754] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1960 < i_size && h_count >= i_worm_x[11765:11760] * PIXEL_SIZE && h_count < i_worm_x[11765:11760] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11765:11760] * PIXEL_SIZE && v_count < i_worm_y[11765:11760] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1961 < i_size && h_count >= i_worm_x[11771:11766] * PIXEL_SIZE && h_count < i_worm_x[11771:11766] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11771:11766] * PIXEL_SIZE && v_count < i_worm_y[11771:11766] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1962 < i_size && h_count >= i_worm_x[11777:11772] * PIXEL_SIZE && h_count < i_worm_x[11777:11772] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11777:11772] * PIXEL_SIZE && v_count < i_worm_y[11777:11772] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1963 < i_size && h_count >= i_worm_x[11783:11778] * PIXEL_SIZE && h_count < i_worm_x[11783:11778] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11783:11778] * PIXEL_SIZE && v_count < i_worm_y[11783:11778] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1964 < i_size && h_count >= i_worm_x[11789:11784] * PIXEL_SIZE && h_count < i_worm_x[11789:11784] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11789:11784] * PIXEL_SIZE && v_count < i_worm_y[11789:11784] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1965 < i_size && h_count >= i_worm_x[11795:11790] * PIXEL_SIZE && h_count < i_worm_x[11795:11790] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11795:11790] * PIXEL_SIZE && v_count < i_worm_y[11795:11790] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1966 < i_size && h_count >= i_worm_x[11801:11796] * PIXEL_SIZE && h_count < i_worm_x[11801:11796] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11801:11796] * PIXEL_SIZE && v_count < i_worm_y[11801:11796] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1967 < i_size && h_count >= i_worm_x[11807:11802] * PIXEL_SIZE && h_count < i_worm_x[11807:11802] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11807:11802] * PIXEL_SIZE && v_count < i_worm_y[11807:11802] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1968 < i_size && h_count >= i_worm_x[11813:11808] * PIXEL_SIZE && h_count < i_worm_x[11813:11808] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11813:11808] * PIXEL_SIZE && v_count < i_worm_y[11813:11808] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1969 < i_size && h_count >= i_worm_x[11819:11814] * PIXEL_SIZE && h_count < i_worm_x[11819:11814] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11819:11814] * PIXEL_SIZE && v_count < i_worm_y[11819:11814] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1970 < i_size && h_count >= i_worm_x[11825:11820] * PIXEL_SIZE && h_count < i_worm_x[11825:11820] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11825:11820] * PIXEL_SIZE && v_count < i_worm_y[11825:11820] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1971 < i_size && h_count >= i_worm_x[11831:11826] * PIXEL_SIZE && h_count < i_worm_x[11831:11826] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11831:11826] * PIXEL_SIZE && v_count < i_worm_y[11831:11826] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1972 < i_size && h_count >= i_worm_x[11837:11832] * PIXEL_SIZE && h_count < i_worm_x[11837:11832] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11837:11832] * PIXEL_SIZE && v_count < i_worm_y[11837:11832] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1973 < i_size && h_count >= i_worm_x[11843:11838] * PIXEL_SIZE && h_count < i_worm_x[11843:11838] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11843:11838] * PIXEL_SIZE && v_count < i_worm_y[11843:11838] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1974 < i_size && h_count >= i_worm_x[11849:11844] * PIXEL_SIZE && h_count < i_worm_x[11849:11844] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11849:11844] * PIXEL_SIZE && v_count < i_worm_y[11849:11844] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1975 < i_size && h_count >= i_worm_x[11855:11850] * PIXEL_SIZE && h_count < i_worm_x[11855:11850] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11855:11850] * PIXEL_SIZE && v_count < i_worm_y[11855:11850] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1976 < i_size && h_count >= i_worm_x[11861:11856] * PIXEL_SIZE && h_count < i_worm_x[11861:11856] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11861:11856] * PIXEL_SIZE && v_count < i_worm_y[11861:11856] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1977 < i_size && h_count >= i_worm_x[11867:11862] * PIXEL_SIZE && h_count < i_worm_x[11867:11862] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11867:11862] * PIXEL_SIZE && v_count < i_worm_y[11867:11862] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1978 < i_size && h_count >= i_worm_x[11873:11868] * PIXEL_SIZE && h_count < i_worm_x[11873:11868] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11873:11868] * PIXEL_SIZE && v_count < i_worm_y[11873:11868] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1979 < i_size && h_count >= i_worm_x[11879:11874] * PIXEL_SIZE && h_count < i_worm_x[11879:11874] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11879:11874] * PIXEL_SIZE && v_count < i_worm_y[11879:11874] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1980 < i_size && h_count >= i_worm_x[11885:11880] * PIXEL_SIZE && h_count < i_worm_x[11885:11880] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11885:11880] * PIXEL_SIZE && v_count < i_worm_y[11885:11880] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1981 < i_size && h_count >= i_worm_x[11891:11886] * PIXEL_SIZE && h_count < i_worm_x[11891:11886] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11891:11886] * PIXEL_SIZE && v_count < i_worm_y[11891:11886] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1982 < i_size && h_count >= i_worm_x[11897:11892] * PIXEL_SIZE && h_count < i_worm_x[11897:11892] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11897:11892] * PIXEL_SIZE && v_count < i_worm_y[11897:11892] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1983 < i_size && h_count >= i_worm_x[11903:11898] * PIXEL_SIZE && h_count < i_worm_x[11903:11898] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11903:11898] * PIXEL_SIZE && v_count < i_worm_y[11903:11898] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1984 < i_size && h_count >= i_worm_x[11909:11904] * PIXEL_SIZE && h_count < i_worm_x[11909:11904] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11909:11904] * PIXEL_SIZE && v_count < i_worm_y[11909:11904] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1985 < i_size && h_count >= i_worm_x[11915:11910] * PIXEL_SIZE && h_count < i_worm_x[11915:11910] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11915:11910] * PIXEL_SIZE && v_count < i_worm_y[11915:11910] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1986 < i_size && h_count >= i_worm_x[11921:11916] * PIXEL_SIZE && h_count < i_worm_x[11921:11916] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11921:11916] * PIXEL_SIZE && v_count < i_worm_y[11921:11916] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1987 < i_size && h_count >= i_worm_x[11927:11922] * PIXEL_SIZE && h_count < i_worm_x[11927:11922] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11927:11922] * PIXEL_SIZE && v_count < i_worm_y[11927:11922] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1988 < i_size && h_count >= i_worm_x[11933:11928] * PIXEL_SIZE && h_count < i_worm_x[11933:11928] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11933:11928] * PIXEL_SIZE && v_count < i_worm_y[11933:11928] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1989 < i_size && h_count >= i_worm_x[11939:11934] * PIXEL_SIZE && h_count < i_worm_x[11939:11934] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11939:11934] * PIXEL_SIZE && v_count < i_worm_y[11939:11934] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1990 < i_size && h_count >= i_worm_x[11945:11940] * PIXEL_SIZE && h_count < i_worm_x[11945:11940] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11945:11940] * PIXEL_SIZE && v_count < i_worm_y[11945:11940] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1991 < i_size && h_count >= i_worm_x[11951:11946] * PIXEL_SIZE && h_count < i_worm_x[11951:11946] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11951:11946] * PIXEL_SIZE && v_count < i_worm_y[11951:11946] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1992 < i_size && h_count >= i_worm_x[11957:11952] * PIXEL_SIZE && h_count < i_worm_x[11957:11952] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11957:11952] * PIXEL_SIZE && v_count < i_worm_y[11957:11952] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1993 < i_size && h_count >= i_worm_x[11963:11958] * PIXEL_SIZE && h_count < i_worm_x[11963:11958] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11963:11958] * PIXEL_SIZE && v_count < i_worm_y[11963:11958] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1994 < i_size && h_count >= i_worm_x[11969:11964] * PIXEL_SIZE && h_count < i_worm_x[11969:11964] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11969:11964] * PIXEL_SIZE && v_count < i_worm_y[11969:11964] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1995 < i_size && h_count >= i_worm_x[11975:11970] * PIXEL_SIZE && h_count < i_worm_x[11975:11970] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11975:11970] * PIXEL_SIZE && v_count < i_worm_y[11975:11970] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1996 < i_size && h_count >= i_worm_x[11981:11976] * PIXEL_SIZE && h_count < i_worm_x[11981:11976] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11981:11976] * PIXEL_SIZE && v_count < i_worm_y[11981:11976] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1997 < i_size && h_count >= i_worm_x[11987:11982] * PIXEL_SIZE && h_count < i_worm_x[11987:11982] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11987:11982] * PIXEL_SIZE && v_count < i_worm_y[11987:11982] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1998 < i_size && h_count >= i_worm_x[11993:11988] * PIXEL_SIZE && h_count < i_worm_x[11993:11988] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11993:11988] * PIXEL_SIZE && v_count < i_worm_y[11993:11988] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (1999 < i_size && h_count >= i_worm_x[11999:11994] * PIXEL_SIZE && h_count < i_worm_x[11999:11994] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[11999:11994] * PIXEL_SIZE && v_count < i_worm_y[11999:11994] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2000 < i_size && h_count >= i_worm_x[12005:12000] * PIXEL_SIZE && h_count < i_worm_x[12005:12000] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12005:12000] * PIXEL_SIZE && v_count < i_worm_y[12005:12000] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2001 < i_size && h_count >= i_worm_x[12011:12006] * PIXEL_SIZE && h_count < i_worm_x[12011:12006] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12011:12006] * PIXEL_SIZE && v_count < i_worm_y[12011:12006] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2002 < i_size && h_count >= i_worm_x[12017:12012] * PIXEL_SIZE && h_count < i_worm_x[12017:12012] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12017:12012] * PIXEL_SIZE && v_count < i_worm_y[12017:12012] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2003 < i_size && h_count >= i_worm_x[12023:12018] * PIXEL_SIZE && h_count < i_worm_x[12023:12018] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12023:12018] * PIXEL_SIZE && v_count < i_worm_y[12023:12018] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2004 < i_size && h_count >= i_worm_x[12029:12024] * PIXEL_SIZE && h_count < i_worm_x[12029:12024] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12029:12024] * PIXEL_SIZE && v_count < i_worm_y[12029:12024] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2005 < i_size && h_count >= i_worm_x[12035:12030] * PIXEL_SIZE && h_count < i_worm_x[12035:12030] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12035:12030] * PIXEL_SIZE && v_count < i_worm_y[12035:12030] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2006 < i_size && h_count >= i_worm_x[12041:12036] * PIXEL_SIZE && h_count < i_worm_x[12041:12036] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12041:12036] * PIXEL_SIZE && v_count < i_worm_y[12041:12036] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2007 < i_size && h_count >= i_worm_x[12047:12042] * PIXEL_SIZE && h_count < i_worm_x[12047:12042] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12047:12042] * PIXEL_SIZE && v_count < i_worm_y[12047:12042] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2008 < i_size && h_count >= i_worm_x[12053:12048] * PIXEL_SIZE && h_count < i_worm_x[12053:12048] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12053:12048] * PIXEL_SIZE && v_count < i_worm_y[12053:12048] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2009 < i_size && h_count >= i_worm_x[12059:12054] * PIXEL_SIZE && h_count < i_worm_x[12059:12054] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12059:12054] * PIXEL_SIZE && v_count < i_worm_y[12059:12054] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2010 < i_size && h_count >= i_worm_x[12065:12060] * PIXEL_SIZE && h_count < i_worm_x[12065:12060] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12065:12060] * PIXEL_SIZE && v_count < i_worm_y[12065:12060] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2011 < i_size && h_count >= i_worm_x[12071:12066] * PIXEL_SIZE && h_count < i_worm_x[12071:12066] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12071:12066] * PIXEL_SIZE && v_count < i_worm_y[12071:12066] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2012 < i_size && h_count >= i_worm_x[12077:12072] * PIXEL_SIZE && h_count < i_worm_x[12077:12072] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12077:12072] * PIXEL_SIZE && v_count < i_worm_y[12077:12072] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2013 < i_size && h_count >= i_worm_x[12083:12078] * PIXEL_SIZE && h_count < i_worm_x[12083:12078] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12083:12078] * PIXEL_SIZE && v_count < i_worm_y[12083:12078] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2014 < i_size && h_count >= i_worm_x[12089:12084] * PIXEL_SIZE && h_count < i_worm_x[12089:12084] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12089:12084] * PIXEL_SIZE && v_count < i_worm_y[12089:12084] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2015 < i_size && h_count >= i_worm_x[12095:12090] * PIXEL_SIZE && h_count < i_worm_x[12095:12090] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12095:12090] * PIXEL_SIZE && v_count < i_worm_y[12095:12090] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2016 < i_size && h_count >= i_worm_x[12101:12096] * PIXEL_SIZE && h_count < i_worm_x[12101:12096] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12101:12096] * PIXEL_SIZE && v_count < i_worm_y[12101:12096] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2017 < i_size && h_count >= i_worm_x[12107:12102] * PIXEL_SIZE && h_count < i_worm_x[12107:12102] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12107:12102] * PIXEL_SIZE && v_count < i_worm_y[12107:12102] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2018 < i_size && h_count >= i_worm_x[12113:12108] * PIXEL_SIZE && h_count < i_worm_x[12113:12108] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12113:12108] * PIXEL_SIZE && v_count < i_worm_y[12113:12108] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2019 < i_size && h_count >= i_worm_x[12119:12114] * PIXEL_SIZE && h_count < i_worm_x[12119:12114] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12119:12114] * PIXEL_SIZE && v_count < i_worm_y[12119:12114] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2020 < i_size && h_count >= i_worm_x[12125:12120] * PIXEL_SIZE && h_count < i_worm_x[12125:12120] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12125:12120] * PIXEL_SIZE && v_count < i_worm_y[12125:12120] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2021 < i_size && h_count >= i_worm_x[12131:12126] * PIXEL_SIZE && h_count < i_worm_x[12131:12126] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12131:12126] * PIXEL_SIZE && v_count < i_worm_y[12131:12126] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2022 < i_size && h_count >= i_worm_x[12137:12132] * PIXEL_SIZE && h_count < i_worm_x[12137:12132] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12137:12132] * PIXEL_SIZE && v_count < i_worm_y[12137:12132] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2023 < i_size && h_count >= i_worm_x[12143:12138] * PIXEL_SIZE && h_count < i_worm_x[12143:12138] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12143:12138] * PIXEL_SIZE && v_count < i_worm_y[12143:12138] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2024 < i_size && h_count >= i_worm_x[12149:12144] * PIXEL_SIZE && h_count < i_worm_x[12149:12144] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12149:12144] * PIXEL_SIZE && v_count < i_worm_y[12149:12144] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2025 < i_size && h_count >= i_worm_x[12155:12150] * PIXEL_SIZE && h_count < i_worm_x[12155:12150] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12155:12150] * PIXEL_SIZE && v_count < i_worm_y[12155:12150] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2026 < i_size && h_count >= i_worm_x[12161:12156] * PIXEL_SIZE && h_count < i_worm_x[12161:12156] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12161:12156] * PIXEL_SIZE && v_count < i_worm_y[12161:12156] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2027 < i_size && h_count >= i_worm_x[12167:12162] * PIXEL_SIZE && h_count < i_worm_x[12167:12162] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12167:12162] * PIXEL_SIZE && v_count < i_worm_y[12167:12162] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2028 < i_size && h_count >= i_worm_x[12173:12168] * PIXEL_SIZE && h_count < i_worm_x[12173:12168] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12173:12168] * PIXEL_SIZE && v_count < i_worm_y[12173:12168] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2029 < i_size && h_count >= i_worm_x[12179:12174] * PIXEL_SIZE && h_count < i_worm_x[12179:12174] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12179:12174] * PIXEL_SIZE && v_count < i_worm_y[12179:12174] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2030 < i_size && h_count >= i_worm_x[12185:12180] * PIXEL_SIZE && h_count < i_worm_x[12185:12180] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12185:12180] * PIXEL_SIZE && v_count < i_worm_y[12185:12180] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2031 < i_size && h_count >= i_worm_x[12191:12186] * PIXEL_SIZE && h_count < i_worm_x[12191:12186] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12191:12186] * PIXEL_SIZE && v_count < i_worm_y[12191:12186] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2032 < i_size && h_count >= i_worm_x[12197:12192] * PIXEL_SIZE && h_count < i_worm_x[12197:12192] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12197:12192] * PIXEL_SIZE && v_count < i_worm_y[12197:12192] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2033 < i_size && h_count >= i_worm_x[12203:12198] * PIXEL_SIZE && h_count < i_worm_x[12203:12198] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12203:12198] * PIXEL_SIZE && v_count < i_worm_y[12203:12198] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2034 < i_size && h_count >= i_worm_x[12209:12204] * PIXEL_SIZE && h_count < i_worm_x[12209:12204] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12209:12204] * PIXEL_SIZE && v_count < i_worm_y[12209:12204] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2035 < i_size && h_count >= i_worm_x[12215:12210] * PIXEL_SIZE && h_count < i_worm_x[12215:12210] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12215:12210] * PIXEL_SIZE && v_count < i_worm_y[12215:12210] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2036 < i_size && h_count >= i_worm_x[12221:12216] * PIXEL_SIZE && h_count < i_worm_x[12221:12216] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12221:12216] * PIXEL_SIZE && v_count < i_worm_y[12221:12216] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2037 < i_size && h_count >= i_worm_x[12227:12222] * PIXEL_SIZE && h_count < i_worm_x[12227:12222] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12227:12222] * PIXEL_SIZE && v_count < i_worm_y[12227:12222] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2038 < i_size && h_count >= i_worm_x[12233:12228] * PIXEL_SIZE && h_count < i_worm_x[12233:12228] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12233:12228] * PIXEL_SIZE && v_count < i_worm_y[12233:12228] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2039 < i_size && h_count >= i_worm_x[12239:12234] * PIXEL_SIZE && h_count < i_worm_x[12239:12234] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12239:12234] * PIXEL_SIZE && v_count < i_worm_y[12239:12234] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2040 < i_size && h_count >= i_worm_x[12245:12240] * PIXEL_SIZE && h_count < i_worm_x[12245:12240] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12245:12240] * PIXEL_SIZE && v_count < i_worm_y[12245:12240] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2041 < i_size && h_count >= i_worm_x[12251:12246] * PIXEL_SIZE && h_count < i_worm_x[12251:12246] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12251:12246] * PIXEL_SIZE && v_count < i_worm_y[12251:12246] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2042 < i_size && h_count >= i_worm_x[12257:12252] * PIXEL_SIZE && h_count < i_worm_x[12257:12252] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12257:12252] * PIXEL_SIZE && v_count < i_worm_y[12257:12252] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2043 < i_size && h_count >= i_worm_x[12263:12258] * PIXEL_SIZE && h_count < i_worm_x[12263:12258] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12263:12258] * PIXEL_SIZE && v_count < i_worm_y[12263:12258] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2044 < i_size && h_count >= i_worm_x[12269:12264] * PIXEL_SIZE && h_count < i_worm_x[12269:12264] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12269:12264] * PIXEL_SIZE && v_count < i_worm_y[12269:12264] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2045 < i_size && h_count >= i_worm_x[12275:12270] * PIXEL_SIZE && h_count < i_worm_x[12275:12270] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12275:12270] * PIXEL_SIZE && v_count < i_worm_y[12275:12270] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2046 < i_size && h_count >= i_worm_x[12281:12276] * PIXEL_SIZE && h_count < i_worm_x[12281:12276] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12281:12276] * PIXEL_SIZE && v_count < i_worm_y[12281:12276] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2047 < i_size && h_count >= i_worm_x[12287:12282] * PIXEL_SIZE && h_count < i_worm_x[12287:12282] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12287:12282] * PIXEL_SIZE && v_count < i_worm_y[12287:12282] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2048 < i_size && h_count >= i_worm_x[12293:12288] * PIXEL_SIZE && h_count < i_worm_x[12293:12288] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12293:12288] * PIXEL_SIZE && v_count < i_worm_y[12293:12288] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2049 < i_size && h_count >= i_worm_x[12299:12294] * PIXEL_SIZE && h_count < i_worm_x[12299:12294] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12299:12294] * PIXEL_SIZE && v_count < i_worm_y[12299:12294] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2050 < i_size && h_count >= i_worm_x[12305:12300] * PIXEL_SIZE && h_count < i_worm_x[12305:12300] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12305:12300] * PIXEL_SIZE && v_count < i_worm_y[12305:12300] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2051 < i_size && h_count >= i_worm_x[12311:12306] * PIXEL_SIZE && h_count < i_worm_x[12311:12306] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12311:12306] * PIXEL_SIZE && v_count < i_worm_y[12311:12306] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2052 < i_size && h_count >= i_worm_x[12317:12312] * PIXEL_SIZE && h_count < i_worm_x[12317:12312] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12317:12312] * PIXEL_SIZE && v_count < i_worm_y[12317:12312] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2053 < i_size && h_count >= i_worm_x[12323:12318] * PIXEL_SIZE && h_count < i_worm_x[12323:12318] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12323:12318] * PIXEL_SIZE && v_count < i_worm_y[12323:12318] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2054 < i_size && h_count >= i_worm_x[12329:12324] * PIXEL_SIZE && h_count < i_worm_x[12329:12324] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12329:12324] * PIXEL_SIZE && v_count < i_worm_y[12329:12324] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2055 < i_size && h_count >= i_worm_x[12335:12330] * PIXEL_SIZE && h_count < i_worm_x[12335:12330] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12335:12330] * PIXEL_SIZE && v_count < i_worm_y[12335:12330] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2056 < i_size && h_count >= i_worm_x[12341:12336] * PIXEL_SIZE && h_count < i_worm_x[12341:12336] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12341:12336] * PIXEL_SIZE && v_count < i_worm_y[12341:12336] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2057 < i_size && h_count >= i_worm_x[12347:12342] * PIXEL_SIZE && h_count < i_worm_x[12347:12342] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12347:12342] * PIXEL_SIZE && v_count < i_worm_y[12347:12342] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2058 < i_size && h_count >= i_worm_x[12353:12348] * PIXEL_SIZE && h_count < i_worm_x[12353:12348] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12353:12348] * PIXEL_SIZE && v_count < i_worm_y[12353:12348] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2059 < i_size && h_count >= i_worm_x[12359:12354] * PIXEL_SIZE && h_count < i_worm_x[12359:12354] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12359:12354] * PIXEL_SIZE && v_count < i_worm_y[12359:12354] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2060 < i_size && h_count >= i_worm_x[12365:12360] * PIXEL_SIZE && h_count < i_worm_x[12365:12360] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12365:12360] * PIXEL_SIZE && v_count < i_worm_y[12365:12360] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2061 < i_size && h_count >= i_worm_x[12371:12366] * PIXEL_SIZE && h_count < i_worm_x[12371:12366] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12371:12366] * PIXEL_SIZE && v_count < i_worm_y[12371:12366] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2062 < i_size && h_count >= i_worm_x[12377:12372] * PIXEL_SIZE && h_count < i_worm_x[12377:12372] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12377:12372] * PIXEL_SIZE && v_count < i_worm_y[12377:12372] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2063 < i_size && h_count >= i_worm_x[12383:12378] * PIXEL_SIZE && h_count < i_worm_x[12383:12378] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12383:12378] * PIXEL_SIZE && v_count < i_worm_y[12383:12378] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2064 < i_size && h_count >= i_worm_x[12389:12384] * PIXEL_SIZE && h_count < i_worm_x[12389:12384] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12389:12384] * PIXEL_SIZE && v_count < i_worm_y[12389:12384] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2065 < i_size && h_count >= i_worm_x[12395:12390] * PIXEL_SIZE && h_count < i_worm_x[12395:12390] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12395:12390] * PIXEL_SIZE && v_count < i_worm_y[12395:12390] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2066 < i_size && h_count >= i_worm_x[12401:12396] * PIXEL_SIZE && h_count < i_worm_x[12401:12396] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12401:12396] * PIXEL_SIZE && v_count < i_worm_y[12401:12396] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2067 < i_size && h_count >= i_worm_x[12407:12402] * PIXEL_SIZE && h_count < i_worm_x[12407:12402] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12407:12402] * PIXEL_SIZE && v_count < i_worm_y[12407:12402] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2068 < i_size && h_count >= i_worm_x[12413:12408] * PIXEL_SIZE && h_count < i_worm_x[12413:12408] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12413:12408] * PIXEL_SIZE && v_count < i_worm_y[12413:12408] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2069 < i_size && h_count >= i_worm_x[12419:12414] * PIXEL_SIZE && h_count < i_worm_x[12419:12414] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12419:12414] * PIXEL_SIZE && v_count < i_worm_y[12419:12414] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2070 < i_size && h_count >= i_worm_x[12425:12420] * PIXEL_SIZE && h_count < i_worm_x[12425:12420] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12425:12420] * PIXEL_SIZE && v_count < i_worm_y[12425:12420] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2071 < i_size && h_count >= i_worm_x[12431:12426] * PIXEL_SIZE && h_count < i_worm_x[12431:12426] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12431:12426] * PIXEL_SIZE && v_count < i_worm_y[12431:12426] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2072 < i_size && h_count >= i_worm_x[12437:12432] * PIXEL_SIZE && h_count < i_worm_x[12437:12432] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12437:12432] * PIXEL_SIZE && v_count < i_worm_y[12437:12432] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2073 < i_size && h_count >= i_worm_x[12443:12438] * PIXEL_SIZE && h_count < i_worm_x[12443:12438] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12443:12438] * PIXEL_SIZE && v_count < i_worm_y[12443:12438] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2074 < i_size && h_count >= i_worm_x[12449:12444] * PIXEL_SIZE && h_count < i_worm_x[12449:12444] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12449:12444] * PIXEL_SIZE && v_count < i_worm_y[12449:12444] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2075 < i_size && h_count >= i_worm_x[12455:12450] * PIXEL_SIZE && h_count < i_worm_x[12455:12450] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12455:12450] * PIXEL_SIZE && v_count < i_worm_y[12455:12450] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2076 < i_size && h_count >= i_worm_x[12461:12456] * PIXEL_SIZE && h_count < i_worm_x[12461:12456] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12461:12456] * PIXEL_SIZE && v_count < i_worm_y[12461:12456] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2077 < i_size && h_count >= i_worm_x[12467:12462] * PIXEL_SIZE && h_count < i_worm_x[12467:12462] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12467:12462] * PIXEL_SIZE && v_count < i_worm_y[12467:12462] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2078 < i_size && h_count >= i_worm_x[12473:12468] * PIXEL_SIZE && h_count < i_worm_x[12473:12468] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12473:12468] * PIXEL_SIZE && v_count < i_worm_y[12473:12468] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2079 < i_size && h_count >= i_worm_x[12479:12474] * PIXEL_SIZE && h_count < i_worm_x[12479:12474] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12479:12474] * PIXEL_SIZE && v_count < i_worm_y[12479:12474] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2080 < i_size && h_count >= i_worm_x[12485:12480] * PIXEL_SIZE && h_count < i_worm_x[12485:12480] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12485:12480] * PIXEL_SIZE && v_count < i_worm_y[12485:12480] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2081 < i_size && h_count >= i_worm_x[12491:12486] * PIXEL_SIZE && h_count < i_worm_x[12491:12486] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12491:12486] * PIXEL_SIZE && v_count < i_worm_y[12491:12486] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2082 < i_size && h_count >= i_worm_x[12497:12492] * PIXEL_SIZE && h_count < i_worm_x[12497:12492] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12497:12492] * PIXEL_SIZE && v_count < i_worm_y[12497:12492] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2083 < i_size && h_count >= i_worm_x[12503:12498] * PIXEL_SIZE && h_count < i_worm_x[12503:12498] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12503:12498] * PIXEL_SIZE && v_count < i_worm_y[12503:12498] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2084 < i_size && h_count >= i_worm_x[12509:12504] * PIXEL_SIZE && h_count < i_worm_x[12509:12504] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12509:12504] * PIXEL_SIZE && v_count < i_worm_y[12509:12504] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2085 < i_size && h_count >= i_worm_x[12515:12510] * PIXEL_SIZE && h_count < i_worm_x[12515:12510] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12515:12510] * PIXEL_SIZE && v_count < i_worm_y[12515:12510] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2086 < i_size && h_count >= i_worm_x[12521:12516] * PIXEL_SIZE && h_count < i_worm_x[12521:12516] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12521:12516] * PIXEL_SIZE && v_count < i_worm_y[12521:12516] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2087 < i_size && h_count >= i_worm_x[12527:12522] * PIXEL_SIZE && h_count < i_worm_x[12527:12522] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12527:12522] * PIXEL_SIZE && v_count < i_worm_y[12527:12522] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2088 < i_size && h_count >= i_worm_x[12533:12528] * PIXEL_SIZE && h_count < i_worm_x[12533:12528] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12533:12528] * PIXEL_SIZE && v_count < i_worm_y[12533:12528] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2089 < i_size && h_count >= i_worm_x[12539:12534] * PIXEL_SIZE && h_count < i_worm_x[12539:12534] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12539:12534] * PIXEL_SIZE && v_count < i_worm_y[12539:12534] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2090 < i_size && h_count >= i_worm_x[12545:12540] * PIXEL_SIZE && h_count < i_worm_x[12545:12540] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12545:12540] * PIXEL_SIZE && v_count < i_worm_y[12545:12540] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2091 < i_size && h_count >= i_worm_x[12551:12546] * PIXEL_SIZE && h_count < i_worm_x[12551:12546] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12551:12546] * PIXEL_SIZE && v_count < i_worm_y[12551:12546] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2092 < i_size && h_count >= i_worm_x[12557:12552] * PIXEL_SIZE && h_count < i_worm_x[12557:12552] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12557:12552] * PIXEL_SIZE && v_count < i_worm_y[12557:12552] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2093 < i_size && h_count >= i_worm_x[12563:12558] * PIXEL_SIZE && h_count < i_worm_x[12563:12558] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12563:12558] * PIXEL_SIZE && v_count < i_worm_y[12563:12558] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2094 < i_size && h_count >= i_worm_x[12569:12564] * PIXEL_SIZE && h_count < i_worm_x[12569:12564] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12569:12564] * PIXEL_SIZE && v_count < i_worm_y[12569:12564] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2095 < i_size && h_count >= i_worm_x[12575:12570] * PIXEL_SIZE && h_count < i_worm_x[12575:12570] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12575:12570] * PIXEL_SIZE && v_count < i_worm_y[12575:12570] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2096 < i_size && h_count >= i_worm_x[12581:12576] * PIXEL_SIZE && h_count < i_worm_x[12581:12576] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12581:12576] * PIXEL_SIZE && v_count < i_worm_y[12581:12576] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2097 < i_size && h_count >= i_worm_x[12587:12582] * PIXEL_SIZE && h_count < i_worm_x[12587:12582] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12587:12582] * PIXEL_SIZE && v_count < i_worm_y[12587:12582] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2098 < i_size && h_count >= i_worm_x[12593:12588] * PIXEL_SIZE && h_count < i_worm_x[12593:12588] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12593:12588] * PIXEL_SIZE && v_count < i_worm_y[12593:12588] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2099 < i_size && h_count >= i_worm_x[12599:12594] * PIXEL_SIZE && h_count < i_worm_x[12599:12594] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12599:12594] * PIXEL_SIZE && v_count < i_worm_y[12599:12594] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2100 < i_size && h_count >= i_worm_x[12605:12600] * PIXEL_SIZE && h_count < i_worm_x[12605:12600] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12605:12600] * PIXEL_SIZE && v_count < i_worm_y[12605:12600] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2101 < i_size && h_count >= i_worm_x[12611:12606] * PIXEL_SIZE && h_count < i_worm_x[12611:12606] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12611:12606] * PIXEL_SIZE && v_count < i_worm_y[12611:12606] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2102 < i_size && h_count >= i_worm_x[12617:12612] * PIXEL_SIZE && h_count < i_worm_x[12617:12612] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12617:12612] * PIXEL_SIZE && v_count < i_worm_y[12617:12612] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2103 < i_size && h_count >= i_worm_x[12623:12618] * PIXEL_SIZE && h_count < i_worm_x[12623:12618] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12623:12618] * PIXEL_SIZE && v_count < i_worm_y[12623:12618] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2104 < i_size && h_count >= i_worm_x[12629:12624] * PIXEL_SIZE && h_count < i_worm_x[12629:12624] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12629:12624] * PIXEL_SIZE && v_count < i_worm_y[12629:12624] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2105 < i_size && h_count >= i_worm_x[12635:12630] * PIXEL_SIZE && h_count < i_worm_x[12635:12630] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12635:12630] * PIXEL_SIZE && v_count < i_worm_y[12635:12630] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2106 < i_size && h_count >= i_worm_x[12641:12636] * PIXEL_SIZE && h_count < i_worm_x[12641:12636] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12641:12636] * PIXEL_SIZE && v_count < i_worm_y[12641:12636] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2107 < i_size && h_count >= i_worm_x[12647:12642] * PIXEL_SIZE && h_count < i_worm_x[12647:12642] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12647:12642] * PIXEL_SIZE && v_count < i_worm_y[12647:12642] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2108 < i_size && h_count >= i_worm_x[12653:12648] * PIXEL_SIZE && h_count < i_worm_x[12653:12648] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12653:12648] * PIXEL_SIZE && v_count < i_worm_y[12653:12648] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2109 < i_size && h_count >= i_worm_x[12659:12654] * PIXEL_SIZE && h_count < i_worm_x[12659:12654] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12659:12654] * PIXEL_SIZE && v_count < i_worm_y[12659:12654] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2110 < i_size && h_count >= i_worm_x[12665:12660] * PIXEL_SIZE && h_count < i_worm_x[12665:12660] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12665:12660] * PIXEL_SIZE && v_count < i_worm_y[12665:12660] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2111 < i_size && h_count >= i_worm_x[12671:12666] * PIXEL_SIZE && h_count < i_worm_x[12671:12666] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12671:12666] * PIXEL_SIZE && v_count < i_worm_y[12671:12666] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2112 < i_size && h_count >= i_worm_x[12677:12672] * PIXEL_SIZE && h_count < i_worm_x[12677:12672] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12677:12672] * PIXEL_SIZE && v_count < i_worm_y[12677:12672] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2113 < i_size && h_count >= i_worm_x[12683:12678] * PIXEL_SIZE && h_count < i_worm_x[12683:12678] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12683:12678] * PIXEL_SIZE && v_count < i_worm_y[12683:12678] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2114 < i_size && h_count >= i_worm_x[12689:12684] * PIXEL_SIZE && h_count < i_worm_x[12689:12684] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12689:12684] * PIXEL_SIZE && v_count < i_worm_y[12689:12684] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2115 < i_size && h_count >= i_worm_x[12695:12690] * PIXEL_SIZE && h_count < i_worm_x[12695:12690] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12695:12690] * PIXEL_SIZE && v_count < i_worm_y[12695:12690] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2116 < i_size && h_count >= i_worm_x[12701:12696] * PIXEL_SIZE && h_count < i_worm_x[12701:12696] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12701:12696] * PIXEL_SIZE && v_count < i_worm_y[12701:12696] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2117 < i_size && h_count >= i_worm_x[12707:12702] * PIXEL_SIZE && h_count < i_worm_x[12707:12702] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12707:12702] * PIXEL_SIZE && v_count < i_worm_y[12707:12702] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2118 < i_size && h_count >= i_worm_x[12713:12708] * PIXEL_SIZE && h_count < i_worm_x[12713:12708] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12713:12708] * PIXEL_SIZE && v_count < i_worm_y[12713:12708] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2119 < i_size && h_count >= i_worm_x[12719:12714] * PIXEL_SIZE && h_count < i_worm_x[12719:12714] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12719:12714] * PIXEL_SIZE && v_count < i_worm_y[12719:12714] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2120 < i_size && h_count >= i_worm_x[12725:12720] * PIXEL_SIZE && h_count < i_worm_x[12725:12720] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12725:12720] * PIXEL_SIZE && v_count < i_worm_y[12725:12720] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2121 < i_size && h_count >= i_worm_x[12731:12726] * PIXEL_SIZE && h_count < i_worm_x[12731:12726] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12731:12726] * PIXEL_SIZE && v_count < i_worm_y[12731:12726] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2122 < i_size && h_count >= i_worm_x[12737:12732] * PIXEL_SIZE && h_count < i_worm_x[12737:12732] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12737:12732] * PIXEL_SIZE && v_count < i_worm_y[12737:12732] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2123 < i_size && h_count >= i_worm_x[12743:12738] * PIXEL_SIZE && h_count < i_worm_x[12743:12738] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12743:12738] * PIXEL_SIZE && v_count < i_worm_y[12743:12738] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2124 < i_size && h_count >= i_worm_x[12749:12744] * PIXEL_SIZE && h_count < i_worm_x[12749:12744] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12749:12744] * PIXEL_SIZE && v_count < i_worm_y[12749:12744] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2125 < i_size && h_count >= i_worm_x[12755:12750] * PIXEL_SIZE && h_count < i_worm_x[12755:12750] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12755:12750] * PIXEL_SIZE && v_count < i_worm_y[12755:12750] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2126 < i_size && h_count >= i_worm_x[12761:12756] * PIXEL_SIZE && h_count < i_worm_x[12761:12756] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12761:12756] * PIXEL_SIZE && v_count < i_worm_y[12761:12756] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2127 < i_size && h_count >= i_worm_x[12767:12762] * PIXEL_SIZE && h_count < i_worm_x[12767:12762] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12767:12762] * PIXEL_SIZE && v_count < i_worm_y[12767:12762] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2128 < i_size && h_count >= i_worm_x[12773:12768] * PIXEL_SIZE && h_count < i_worm_x[12773:12768] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12773:12768] * PIXEL_SIZE && v_count < i_worm_y[12773:12768] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2129 < i_size && h_count >= i_worm_x[12779:12774] * PIXEL_SIZE && h_count < i_worm_x[12779:12774] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12779:12774] * PIXEL_SIZE && v_count < i_worm_y[12779:12774] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2130 < i_size && h_count >= i_worm_x[12785:12780] * PIXEL_SIZE && h_count < i_worm_x[12785:12780] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12785:12780] * PIXEL_SIZE && v_count < i_worm_y[12785:12780] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2131 < i_size && h_count >= i_worm_x[12791:12786] * PIXEL_SIZE && h_count < i_worm_x[12791:12786] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12791:12786] * PIXEL_SIZE && v_count < i_worm_y[12791:12786] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2132 < i_size && h_count >= i_worm_x[12797:12792] * PIXEL_SIZE && h_count < i_worm_x[12797:12792] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12797:12792] * PIXEL_SIZE && v_count < i_worm_y[12797:12792] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2133 < i_size && h_count >= i_worm_x[12803:12798] * PIXEL_SIZE && h_count < i_worm_x[12803:12798] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12803:12798] * PIXEL_SIZE && v_count < i_worm_y[12803:12798] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2134 < i_size && h_count >= i_worm_x[12809:12804] * PIXEL_SIZE && h_count < i_worm_x[12809:12804] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12809:12804] * PIXEL_SIZE && v_count < i_worm_y[12809:12804] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2135 < i_size && h_count >= i_worm_x[12815:12810] * PIXEL_SIZE && h_count < i_worm_x[12815:12810] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12815:12810] * PIXEL_SIZE && v_count < i_worm_y[12815:12810] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2136 < i_size && h_count >= i_worm_x[12821:12816] * PIXEL_SIZE && h_count < i_worm_x[12821:12816] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12821:12816] * PIXEL_SIZE && v_count < i_worm_y[12821:12816] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2137 < i_size && h_count >= i_worm_x[12827:12822] * PIXEL_SIZE && h_count < i_worm_x[12827:12822] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12827:12822] * PIXEL_SIZE && v_count < i_worm_y[12827:12822] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2138 < i_size && h_count >= i_worm_x[12833:12828] * PIXEL_SIZE && h_count < i_worm_x[12833:12828] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12833:12828] * PIXEL_SIZE && v_count < i_worm_y[12833:12828] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2139 < i_size && h_count >= i_worm_x[12839:12834] * PIXEL_SIZE && h_count < i_worm_x[12839:12834] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12839:12834] * PIXEL_SIZE && v_count < i_worm_y[12839:12834] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2140 < i_size && h_count >= i_worm_x[12845:12840] * PIXEL_SIZE && h_count < i_worm_x[12845:12840] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12845:12840] * PIXEL_SIZE && v_count < i_worm_y[12845:12840] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2141 < i_size && h_count >= i_worm_x[12851:12846] * PIXEL_SIZE && h_count < i_worm_x[12851:12846] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12851:12846] * PIXEL_SIZE && v_count < i_worm_y[12851:12846] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2142 < i_size && h_count >= i_worm_x[12857:12852] * PIXEL_SIZE && h_count < i_worm_x[12857:12852] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12857:12852] * PIXEL_SIZE && v_count < i_worm_y[12857:12852] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2143 < i_size && h_count >= i_worm_x[12863:12858] * PIXEL_SIZE && h_count < i_worm_x[12863:12858] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12863:12858] * PIXEL_SIZE && v_count < i_worm_y[12863:12858] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2144 < i_size && h_count >= i_worm_x[12869:12864] * PIXEL_SIZE && h_count < i_worm_x[12869:12864] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12869:12864] * PIXEL_SIZE && v_count < i_worm_y[12869:12864] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2145 < i_size && h_count >= i_worm_x[12875:12870] * PIXEL_SIZE && h_count < i_worm_x[12875:12870] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12875:12870] * PIXEL_SIZE && v_count < i_worm_y[12875:12870] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2146 < i_size && h_count >= i_worm_x[12881:12876] * PIXEL_SIZE && h_count < i_worm_x[12881:12876] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12881:12876] * PIXEL_SIZE && v_count < i_worm_y[12881:12876] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2147 < i_size && h_count >= i_worm_x[12887:12882] * PIXEL_SIZE && h_count < i_worm_x[12887:12882] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12887:12882] * PIXEL_SIZE && v_count < i_worm_y[12887:12882] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2148 < i_size && h_count >= i_worm_x[12893:12888] * PIXEL_SIZE && h_count < i_worm_x[12893:12888] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12893:12888] * PIXEL_SIZE && v_count < i_worm_y[12893:12888] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2149 < i_size && h_count >= i_worm_x[12899:12894] * PIXEL_SIZE && h_count < i_worm_x[12899:12894] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12899:12894] * PIXEL_SIZE && v_count < i_worm_y[12899:12894] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2150 < i_size && h_count >= i_worm_x[12905:12900] * PIXEL_SIZE && h_count < i_worm_x[12905:12900] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12905:12900] * PIXEL_SIZE && v_count < i_worm_y[12905:12900] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2151 < i_size && h_count >= i_worm_x[12911:12906] * PIXEL_SIZE && h_count < i_worm_x[12911:12906] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12911:12906] * PIXEL_SIZE && v_count < i_worm_y[12911:12906] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2152 < i_size && h_count >= i_worm_x[12917:12912] * PIXEL_SIZE && h_count < i_worm_x[12917:12912] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12917:12912] * PIXEL_SIZE && v_count < i_worm_y[12917:12912] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2153 < i_size && h_count >= i_worm_x[12923:12918] * PIXEL_SIZE && h_count < i_worm_x[12923:12918] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12923:12918] * PIXEL_SIZE && v_count < i_worm_y[12923:12918] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2154 < i_size && h_count >= i_worm_x[12929:12924] * PIXEL_SIZE && h_count < i_worm_x[12929:12924] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12929:12924] * PIXEL_SIZE && v_count < i_worm_y[12929:12924] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2155 < i_size && h_count >= i_worm_x[12935:12930] * PIXEL_SIZE && h_count < i_worm_x[12935:12930] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12935:12930] * PIXEL_SIZE && v_count < i_worm_y[12935:12930] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2156 < i_size && h_count >= i_worm_x[12941:12936] * PIXEL_SIZE && h_count < i_worm_x[12941:12936] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12941:12936] * PIXEL_SIZE && v_count < i_worm_y[12941:12936] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2157 < i_size && h_count >= i_worm_x[12947:12942] * PIXEL_SIZE && h_count < i_worm_x[12947:12942] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12947:12942] * PIXEL_SIZE && v_count < i_worm_y[12947:12942] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2158 < i_size && h_count >= i_worm_x[12953:12948] * PIXEL_SIZE && h_count < i_worm_x[12953:12948] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12953:12948] * PIXEL_SIZE && v_count < i_worm_y[12953:12948] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2159 < i_size && h_count >= i_worm_x[12959:12954] * PIXEL_SIZE && h_count < i_worm_x[12959:12954] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12959:12954] * PIXEL_SIZE && v_count < i_worm_y[12959:12954] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2160 < i_size && h_count >= i_worm_x[12965:12960] * PIXEL_SIZE && h_count < i_worm_x[12965:12960] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12965:12960] * PIXEL_SIZE && v_count < i_worm_y[12965:12960] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2161 < i_size && h_count >= i_worm_x[12971:12966] * PIXEL_SIZE && h_count < i_worm_x[12971:12966] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12971:12966] * PIXEL_SIZE && v_count < i_worm_y[12971:12966] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2162 < i_size && h_count >= i_worm_x[12977:12972] * PIXEL_SIZE && h_count < i_worm_x[12977:12972] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12977:12972] * PIXEL_SIZE && v_count < i_worm_y[12977:12972] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2163 < i_size && h_count >= i_worm_x[12983:12978] * PIXEL_SIZE && h_count < i_worm_x[12983:12978] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12983:12978] * PIXEL_SIZE && v_count < i_worm_y[12983:12978] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2164 < i_size && h_count >= i_worm_x[12989:12984] * PIXEL_SIZE && h_count < i_worm_x[12989:12984] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12989:12984] * PIXEL_SIZE && v_count < i_worm_y[12989:12984] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2165 < i_size && h_count >= i_worm_x[12995:12990] * PIXEL_SIZE && h_count < i_worm_x[12995:12990] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[12995:12990] * PIXEL_SIZE && v_count < i_worm_y[12995:12990] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2166 < i_size && h_count >= i_worm_x[13001:12996] * PIXEL_SIZE && h_count < i_worm_x[13001:12996] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13001:12996] * PIXEL_SIZE && v_count < i_worm_y[13001:12996] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2167 < i_size && h_count >= i_worm_x[13007:13002] * PIXEL_SIZE && h_count < i_worm_x[13007:13002] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13007:13002] * PIXEL_SIZE && v_count < i_worm_y[13007:13002] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2168 < i_size && h_count >= i_worm_x[13013:13008] * PIXEL_SIZE && h_count < i_worm_x[13013:13008] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13013:13008] * PIXEL_SIZE && v_count < i_worm_y[13013:13008] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2169 < i_size && h_count >= i_worm_x[13019:13014] * PIXEL_SIZE && h_count < i_worm_x[13019:13014] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13019:13014] * PIXEL_SIZE && v_count < i_worm_y[13019:13014] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2170 < i_size && h_count >= i_worm_x[13025:13020] * PIXEL_SIZE && h_count < i_worm_x[13025:13020] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13025:13020] * PIXEL_SIZE && v_count < i_worm_y[13025:13020] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2171 < i_size && h_count >= i_worm_x[13031:13026] * PIXEL_SIZE && h_count < i_worm_x[13031:13026] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13031:13026] * PIXEL_SIZE && v_count < i_worm_y[13031:13026] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2172 < i_size && h_count >= i_worm_x[13037:13032] * PIXEL_SIZE && h_count < i_worm_x[13037:13032] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13037:13032] * PIXEL_SIZE && v_count < i_worm_y[13037:13032] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2173 < i_size && h_count >= i_worm_x[13043:13038] * PIXEL_SIZE && h_count < i_worm_x[13043:13038] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13043:13038] * PIXEL_SIZE && v_count < i_worm_y[13043:13038] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2174 < i_size && h_count >= i_worm_x[13049:13044] * PIXEL_SIZE && h_count < i_worm_x[13049:13044] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13049:13044] * PIXEL_SIZE && v_count < i_worm_y[13049:13044] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2175 < i_size && h_count >= i_worm_x[13055:13050] * PIXEL_SIZE && h_count < i_worm_x[13055:13050] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13055:13050] * PIXEL_SIZE && v_count < i_worm_y[13055:13050] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2176 < i_size && h_count >= i_worm_x[13061:13056] * PIXEL_SIZE && h_count < i_worm_x[13061:13056] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13061:13056] * PIXEL_SIZE && v_count < i_worm_y[13061:13056] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2177 < i_size && h_count >= i_worm_x[13067:13062] * PIXEL_SIZE && h_count < i_worm_x[13067:13062] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13067:13062] * PIXEL_SIZE && v_count < i_worm_y[13067:13062] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2178 < i_size && h_count >= i_worm_x[13073:13068] * PIXEL_SIZE && h_count < i_worm_x[13073:13068] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13073:13068] * PIXEL_SIZE && v_count < i_worm_y[13073:13068] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2179 < i_size && h_count >= i_worm_x[13079:13074] * PIXEL_SIZE && h_count < i_worm_x[13079:13074] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13079:13074] * PIXEL_SIZE && v_count < i_worm_y[13079:13074] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2180 < i_size && h_count >= i_worm_x[13085:13080] * PIXEL_SIZE && h_count < i_worm_x[13085:13080] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13085:13080] * PIXEL_SIZE && v_count < i_worm_y[13085:13080] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2181 < i_size && h_count >= i_worm_x[13091:13086] * PIXEL_SIZE && h_count < i_worm_x[13091:13086] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13091:13086] * PIXEL_SIZE && v_count < i_worm_y[13091:13086] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2182 < i_size && h_count >= i_worm_x[13097:13092] * PIXEL_SIZE && h_count < i_worm_x[13097:13092] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13097:13092] * PIXEL_SIZE && v_count < i_worm_y[13097:13092] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2183 < i_size && h_count >= i_worm_x[13103:13098] * PIXEL_SIZE && h_count < i_worm_x[13103:13098] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13103:13098] * PIXEL_SIZE && v_count < i_worm_y[13103:13098] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2184 < i_size && h_count >= i_worm_x[13109:13104] * PIXEL_SIZE && h_count < i_worm_x[13109:13104] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13109:13104] * PIXEL_SIZE && v_count < i_worm_y[13109:13104] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2185 < i_size && h_count >= i_worm_x[13115:13110] * PIXEL_SIZE && h_count < i_worm_x[13115:13110] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13115:13110] * PIXEL_SIZE && v_count < i_worm_y[13115:13110] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2186 < i_size && h_count >= i_worm_x[13121:13116] * PIXEL_SIZE && h_count < i_worm_x[13121:13116] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13121:13116] * PIXEL_SIZE && v_count < i_worm_y[13121:13116] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2187 < i_size && h_count >= i_worm_x[13127:13122] * PIXEL_SIZE && h_count < i_worm_x[13127:13122] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13127:13122] * PIXEL_SIZE && v_count < i_worm_y[13127:13122] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2188 < i_size && h_count >= i_worm_x[13133:13128] * PIXEL_SIZE && h_count < i_worm_x[13133:13128] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13133:13128] * PIXEL_SIZE && v_count < i_worm_y[13133:13128] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2189 < i_size && h_count >= i_worm_x[13139:13134] * PIXEL_SIZE && h_count < i_worm_x[13139:13134] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13139:13134] * PIXEL_SIZE && v_count < i_worm_y[13139:13134] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2190 < i_size && h_count >= i_worm_x[13145:13140] * PIXEL_SIZE && h_count < i_worm_x[13145:13140] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13145:13140] * PIXEL_SIZE && v_count < i_worm_y[13145:13140] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2191 < i_size && h_count >= i_worm_x[13151:13146] * PIXEL_SIZE && h_count < i_worm_x[13151:13146] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13151:13146] * PIXEL_SIZE && v_count < i_worm_y[13151:13146] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2192 < i_size && h_count >= i_worm_x[13157:13152] * PIXEL_SIZE && h_count < i_worm_x[13157:13152] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13157:13152] * PIXEL_SIZE && v_count < i_worm_y[13157:13152] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2193 < i_size && h_count >= i_worm_x[13163:13158] * PIXEL_SIZE && h_count < i_worm_x[13163:13158] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13163:13158] * PIXEL_SIZE && v_count < i_worm_y[13163:13158] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2194 < i_size && h_count >= i_worm_x[13169:13164] * PIXEL_SIZE && h_count < i_worm_x[13169:13164] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13169:13164] * PIXEL_SIZE && v_count < i_worm_y[13169:13164] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2195 < i_size && h_count >= i_worm_x[13175:13170] * PIXEL_SIZE && h_count < i_worm_x[13175:13170] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13175:13170] * PIXEL_SIZE && v_count < i_worm_y[13175:13170] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2196 < i_size && h_count >= i_worm_x[13181:13176] * PIXEL_SIZE && h_count < i_worm_x[13181:13176] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13181:13176] * PIXEL_SIZE && v_count < i_worm_y[13181:13176] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2197 < i_size && h_count >= i_worm_x[13187:13182] * PIXEL_SIZE && h_count < i_worm_x[13187:13182] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13187:13182] * PIXEL_SIZE && v_count < i_worm_y[13187:13182] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2198 < i_size && h_count >= i_worm_x[13193:13188] * PIXEL_SIZE && h_count < i_worm_x[13193:13188] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13193:13188] * PIXEL_SIZE && v_count < i_worm_y[13193:13188] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2199 < i_size && h_count >= i_worm_x[13199:13194] * PIXEL_SIZE && h_count < i_worm_x[13199:13194] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13199:13194] * PIXEL_SIZE && v_count < i_worm_y[13199:13194] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2200 < i_size && h_count >= i_worm_x[13205:13200] * PIXEL_SIZE && h_count < i_worm_x[13205:13200] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13205:13200] * PIXEL_SIZE && v_count < i_worm_y[13205:13200] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2201 < i_size && h_count >= i_worm_x[13211:13206] * PIXEL_SIZE && h_count < i_worm_x[13211:13206] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13211:13206] * PIXEL_SIZE && v_count < i_worm_y[13211:13206] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2202 < i_size && h_count >= i_worm_x[13217:13212] * PIXEL_SIZE && h_count < i_worm_x[13217:13212] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13217:13212] * PIXEL_SIZE && v_count < i_worm_y[13217:13212] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2203 < i_size && h_count >= i_worm_x[13223:13218] * PIXEL_SIZE && h_count < i_worm_x[13223:13218] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13223:13218] * PIXEL_SIZE && v_count < i_worm_y[13223:13218] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2204 < i_size && h_count >= i_worm_x[13229:13224] * PIXEL_SIZE && h_count < i_worm_x[13229:13224] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13229:13224] * PIXEL_SIZE && v_count < i_worm_y[13229:13224] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2205 < i_size && h_count >= i_worm_x[13235:13230] * PIXEL_SIZE && h_count < i_worm_x[13235:13230] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13235:13230] * PIXEL_SIZE && v_count < i_worm_y[13235:13230] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2206 < i_size && h_count >= i_worm_x[13241:13236] * PIXEL_SIZE && h_count < i_worm_x[13241:13236] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13241:13236] * PIXEL_SIZE && v_count < i_worm_y[13241:13236] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2207 < i_size && h_count >= i_worm_x[13247:13242] * PIXEL_SIZE && h_count < i_worm_x[13247:13242] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13247:13242] * PIXEL_SIZE && v_count < i_worm_y[13247:13242] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2208 < i_size && h_count >= i_worm_x[13253:13248] * PIXEL_SIZE && h_count < i_worm_x[13253:13248] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13253:13248] * PIXEL_SIZE && v_count < i_worm_y[13253:13248] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2209 < i_size && h_count >= i_worm_x[13259:13254] * PIXEL_SIZE && h_count < i_worm_x[13259:13254] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13259:13254] * PIXEL_SIZE && v_count < i_worm_y[13259:13254] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2210 < i_size && h_count >= i_worm_x[13265:13260] * PIXEL_SIZE && h_count < i_worm_x[13265:13260] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13265:13260] * PIXEL_SIZE && v_count < i_worm_y[13265:13260] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2211 < i_size && h_count >= i_worm_x[13271:13266] * PIXEL_SIZE && h_count < i_worm_x[13271:13266] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13271:13266] * PIXEL_SIZE && v_count < i_worm_y[13271:13266] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2212 < i_size && h_count >= i_worm_x[13277:13272] * PIXEL_SIZE && h_count < i_worm_x[13277:13272] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13277:13272] * PIXEL_SIZE && v_count < i_worm_y[13277:13272] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2213 < i_size && h_count >= i_worm_x[13283:13278] * PIXEL_SIZE && h_count < i_worm_x[13283:13278] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13283:13278] * PIXEL_SIZE && v_count < i_worm_y[13283:13278] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2214 < i_size && h_count >= i_worm_x[13289:13284] * PIXEL_SIZE && h_count < i_worm_x[13289:13284] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13289:13284] * PIXEL_SIZE && v_count < i_worm_y[13289:13284] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2215 < i_size && h_count >= i_worm_x[13295:13290] * PIXEL_SIZE && h_count < i_worm_x[13295:13290] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13295:13290] * PIXEL_SIZE && v_count < i_worm_y[13295:13290] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2216 < i_size && h_count >= i_worm_x[13301:13296] * PIXEL_SIZE && h_count < i_worm_x[13301:13296] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13301:13296] * PIXEL_SIZE && v_count < i_worm_y[13301:13296] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2217 < i_size && h_count >= i_worm_x[13307:13302] * PIXEL_SIZE && h_count < i_worm_x[13307:13302] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13307:13302] * PIXEL_SIZE && v_count < i_worm_y[13307:13302] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2218 < i_size && h_count >= i_worm_x[13313:13308] * PIXEL_SIZE && h_count < i_worm_x[13313:13308] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13313:13308] * PIXEL_SIZE && v_count < i_worm_y[13313:13308] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2219 < i_size && h_count >= i_worm_x[13319:13314] * PIXEL_SIZE && h_count < i_worm_x[13319:13314] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13319:13314] * PIXEL_SIZE && v_count < i_worm_y[13319:13314] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2220 < i_size && h_count >= i_worm_x[13325:13320] * PIXEL_SIZE && h_count < i_worm_x[13325:13320] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13325:13320] * PIXEL_SIZE && v_count < i_worm_y[13325:13320] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2221 < i_size && h_count >= i_worm_x[13331:13326] * PIXEL_SIZE && h_count < i_worm_x[13331:13326] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13331:13326] * PIXEL_SIZE && v_count < i_worm_y[13331:13326] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2222 < i_size && h_count >= i_worm_x[13337:13332] * PIXEL_SIZE && h_count < i_worm_x[13337:13332] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13337:13332] * PIXEL_SIZE && v_count < i_worm_y[13337:13332] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2223 < i_size && h_count >= i_worm_x[13343:13338] * PIXEL_SIZE && h_count < i_worm_x[13343:13338] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13343:13338] * PIXEL_SIZE && v_count < i_worm_y[13343:13338] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2224 < i_size && h_count >= i_worm_x[13349:13344] * PIXEL_SIZE && h_count < i_worm_x[13349:13344] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13349:13344] * PIXEL_SIZE && v_count < i_worm_y[13349:13344] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2225 < i_size && h_count >= i_worm_x[13355:13350] * PIXEL_SIZE && h_count < i_worm_x[13355:13350] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13355:13350] * PIXEL_SIZE && v_count < i_worm_y[13355:13350] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2226 < i_size && h_count >= i_worm_x[13361:13356] * PIXEL_SIZE && h_count < i_worm_x[13361:13356] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13361:13356] * PIXEL_SIZE && v_count < i_worm_y[13361:13356] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2227 < i_size && h_count >= i_worm_x[13367:13362] * PIXEL_SIZE && h_count < i_worm_x[13367:13362] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13367:13362] * PIXEL_SIZE && v_count < i_worm_y[13367:13362] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2228 < i_size && h_count >= i_worm_x[13373:13368] * PIXEL_SIZE && h_count < i_worm_x[13373:13368] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13373:13368] * PIXEL_SIZE && v_count < i_worm_y[13373:13368] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2229 < i_size && h_count >= i_worm_x[13379:13374] * PIXEL_SIZE && h_count < i_worm_x[13379:13374] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13379:13374] * PIXEL_SIZE && v_count < i_worm_y[13379:13374] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2230 < i_size && h_count >= i_worm_x[13385:13380] * PIXEL_SIZE && h_count < i_worm_x[13385:13380] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13385:13380] * PIXEL_SIZE && v_count < i_worm_y[13385:13380] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2231 < i_size && h_count >= i_worm_x[13391:13386] * PIXEL_SIZE && h_count < i_worm_x[13391:13386] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13391:13386] * PIXEL_SIZE && v_count < i_worm_y[13391:13386] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2232 < i_size && h_count >= i_worm_x[13397:13392] * PIXEL_SIZE && h_count < i_worm_x[13397:13392] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13397:13392] * PIXEL_SIZE && v_count < i_worm_y[13397:13392] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2233 < i_size && h_count >= i_worm_x[13403:13398] * PIXEL_SIZE && h_count < i_worm_x[13403:13398] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13403:13398] * PIXEL_SIZE && v_count < i_worm_y[13403:13398] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2234 < i_size && h_count >= i_worm_x[13409:13404] * PIXEL_SIZE && h_count < i_worm_x[13409:13404] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13409:13404] * PIXEL_SIZE && v_count < i_worm_y[13409:13404] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2235 < i_size && h_count >= i_worm_x[13415:13410] * PIXEL_SIZE && h_count < i_worm_x[13415:13410] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13415:13410] * PIXEL_SIZE && v_count < i_worm_y[13415:13410] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2236 < i_size && h_count >= i_worm_x[13421:13416] * PIXEL_SIZE && h_count < i_worm_x[13421:13416] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13421:13416] * PIXEL_SIZE && v_count < i_worm_y[13421:13416] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2237 < i_size && h_count >= i_worm_x[13427:13422] * PIXEL_SIZE && h_count < i_worm_x[13427:13422] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13427:13422] * PIXEL_SIZE && v_count < i_worm_y[13427:13422] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2238 < i_size && h_count >= i_worm_x[13433:13428] * PIXEL_SIZE && h_count < i_worm_x[13433:13428] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13433:13428] * PIXEL_SIZE && v_count < i_worm_y[13433:13428] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2239 < i_size && h_count >= i_worm_x[13439:13434] * PIXEL_SIZE && h_count < i_worm_x[13439:13434] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13439:13434] * PIXEL_SIZE && v_count < i_worm_y[13439:13434] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2240 < i_size && h_count >= i_worm_x[13445:13440] * PIXEL_SIZE && h_count < i_worm_x[13445:13440] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13445:13440] * PIXEL_SIZE && v_count < i_worm_y[13445:13440] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2241 < i_size && h_count >= i_worm_x[13451:13446] * PIXEL_SIZE && h_count < i_worm_x[13451:13446] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13451:13446] * PIXEL_SIZE && v_count < i_worm_y[13451:13446] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2242 < i_size && h_count >= i_worm_x[13457:13452] * PIXEL_SIZE && h_count < i_worm_x[13457:13452] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13457:13452] * PIXEL_SIZE && v_count < i_worm_y[13457:13452] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2243 < i_size && h_count >= i_worm_x[13463:13458] * PIXEL_SIZE && h_count < i_worm_x[13463:13458] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13463:13458] * PIXEL_SIZE && v_count < i_worm_y[13463:13458] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2244 < i_size && h_count >= i_worm_x[13469:13464] * PIXEL_SIZE && h_count < i_worm_x[13469:13464] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13469:13464] * PIXEL_SIZE && v_count < i_worm_y[13469:13464] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2245 < i_size && h_count >= i_worm_x[13475:13470] * PIXEL_SIZE && h_count < i_worm_x[13475:13470] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13475:13470] * PIXEL_SIZE && v_count < i_worm_y[13475:13470] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2246 < i_size && h_count >= i_worm_x[13481:13476] * PIXEL_SIZE && h_count < i_worm_x[13481:13476] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13481:13476] * PIXEL_SIZE && v_count < i_worm_y[13481:13476] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2247 < i_size && h_count >= i_worm_x[13487:13482] * PIXEL_SIZE && h_count < i_worm_x[13487:13482] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13487:13482] * PIXEL_SIZE && v_count < i_worm_y[13487:13482] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2248 < i_size && h_count >= i_worm_x[13493:13488] * PIXEL_SIZE && h_count < i_worm_x[13493:13488] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13493:13488] * PIXEL_SIZE && v_count < i_worm_y[13493:13488] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2249 < i_size && h_count >= i_worm_x[13499:13494] * PIXEL_SIZE && h_count < i_worm_x[13499:13494] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13499:13494] * PIXEL_SIZE && v_count < i_worm_y[13499:13494] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2250 < i_size && h_count >= i_worm_x[13505:13500] * PIXEL_SIZE && h_count < i_worm_x[13505:13500] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13505:13500] * PIXEL_SIZE && v_count < i_worm_y[13505:13500] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2251 < i_size && h_count >= i_worm_x[13511:13506] * PIXEL_SIZE && h_count < i_worm_x[13511:13506] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13511:13506] * PIXEL_SIZE && v_count < i_worm_y[13511:13506] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2252 < i_size && h_count >= i_worm_x[13517:13512] * PIXEL_SIZE && h_count < i_worm_x[13517:13512] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13517:13512] * PIXEL_SIZE && v_count < i_worm_y[13517:13512] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2253 < i_size && h_count >= i_worm_x[13523:13518] * PIXEL_SIZE && h_count < i_worm_x[13523:13518] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13523:13518] * PIXEL_SIZE && v_count < i_worm_y[13523:13518] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2254 < i_size && h_count >= i_worm_x[13529:13524] * PIXEL_SIZE && h_count < i_worm_x[13529:13524] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13529:13524] * PIXEL_SIZE && v_count < i_worm_y[13529:13524] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2255 < i_size && h_count >= i_worm_x[13535:13530] * PIXEL_SIZE && h_count < i_worm_x[13535:13530] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13535:13530] * PIXEL_SIZE && v_count < i_worm_y[13535:13530] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2256 < i_size && h_count >= i_worm_x[13541:13536] * PIXEL_SIZE && h_count < i_worm_x[13541:13536] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13541:13536] * PIXEL_SIZE && v_count < i_worm_y[13541:13536] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2257 < i_size && h_count >= i_worm_x[13547:13542] * PIXEL_SIZE && h_count < i_worm_x[13547:13542] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13547:13542] * PIXEL_SIZE && v_count < i_worm_y[13547:13542] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2258 < i_size && h_count >= i_worm_x[13553:13548] * PIXEL_SIZE && h_count < i_worm_x[13553:13548] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13553:13548] * PIXEL_SIZE && v_count < i_worm_y[13553:13548] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2259 < i_size && h_count >= i_worm_x[13559:13554] * PIXEL_SIZE && h_count < i_worm_x[13559:13554] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13559:13554] * PIXEL_SIZE && v_count < i_worm_y[13559:13554] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2260 < i_size && h_count >= i_worm_x[13565:13560] * PIXEL_SIZE && h_count < i_worm_x[13565:13560] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13565:13560] * PIXEL_SIZE && v_count < i_worm_y[13565:13560] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2261 < i_size && h_count >= i_worm_x[13571:13566] * PIXEL_SIZE && h_count < i_worm_x[13571:13566] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13571:13566] * PIXEL_SIZE && v_count < i_worm_y[13571:13566] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2262 < i_size && h_count >= i_worm_x[13577:13572] * PIXEL_SIZE && h_count < i_worm_x[13577:13572] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13577:13572] * PIXEL_SIZE && v_count < i_worm_y[13577:13572] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2263 < i_size && h_count >= i_worm_x[13583:13578] * PIXEL_SIZE && h_count < i_worm_x[13583:13578] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13583:13578] * PIXEL_SIZE && v_count < i_worm_y[13583:13578] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2264 < i_size && h_count >= i_worm_x[13589:13584] * PIXEL_SIZE && h_count < i_worm_x[13589:13584] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13589:13584] * PIXEL_SIZE && v_count < i_worm_y[13589:13584] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2265 < i_size && h_count >= i_worm_x[13595:13590] * PIXEL_SIZE && h_count < i_worm_x[13595:13590] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13595:13590] * PIXEL_SIZE && v_count < i_worm_y[13595:13590] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2266 < i_size && h_count >= i_worm_x[13601:13596] * PIXEL_SIZE && h_count < i_worm_x[13601:13596] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13601:13596] * PIXEL_SIZE && v_count < i_worm_y[13601:13596] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2267 < i_size && h_count >= i_worm_x[13607:13602] * PIXEL_SIZE && h_count < i_worm_x[13607:13602] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13607:13602] * PIXEL_SIZE && v_count < i_worm_y[13607:13602] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2268 < i_size && h_count >= i_worm_x[13613:13608] * PIXEL_SIZE && h_count < i_worm_x[13613:13608] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13613:13608] * PIXEL_SIZE && v_count < i_worm_y[13613:13608] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2269 < i_size && h_count >= i_worm_x[13619:13614] * PIXEL_SIZE && h_count < i_worm_x[13619:13614] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13619:13614] * PIXEL_SIZE && v_count < i_worm_y[13619:13614] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2270 < i_size && h_count >= i_worm_x[13625:13620] * PIXEL_SIZE && h_count < i_worm_x[13625:13620] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13625:13620] * PIXEL_SIZE && v_count < i_worm_y[13625:13620] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2271 < i_size && h_count >= i_worm_x[13631:13626] * PIXEL_SIZE && h_count < i_worm_x[13631:13626] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13631:13626] * PIXEL_SIZE && v_count < i_worm_y[13631:13626] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2272 < i_size && h_count >= i_worm_x[13637:13632] * PIXEL_SIZE && h_count < i_worm_x[13637:13632] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13637:13632] * PIXEL_SIZE && v_count < i_worm_y[13637:13632] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2273 < i_size && h_count >= i_worm_x[13643:13638] * PIXEL_SIZE && h_count < i_worm_x[13643:13638] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13643:13638] * PIXEL_SIZE && v_count < i_worm_y[13643:13638] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2274 < i_size && h_count >= i_worm_x[13649:13644] * PIXEL_SIZE && h_count < i_worm_x[13649:13644] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13649:13644] * PIXEL_SIZE && v_count < i_worm_y[13649:13644] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2275 < i_size && h_count >= i_worm_x[13655:13650] * PIXEL_SIZE && h_count < i_worm_x[13655:13650] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13655:13650] * PIXEL_SIZE && v_count < i_worm_y[13655:13650] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2276 < i_size && h_count >= i_worm_x[13661:13656] * PIXEL_SIZE && h_count < i_worm_x[13661:13656] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13661:13656] * PIXEL_SIZE && v_count < i_worm_y[13661:13656] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2277 < i_size && h_count >= i_worm_x[13667:13662] * PIXEL_SIZE && h_count < i_worm_x[13667:13662] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13667:13662] * PIXEL_SIZE && v_count < i_worm_y[13667:13662] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2278 < i_size && h_count >= i_worm_x[13673:13668] * PIXEL_SIZE && h_count < i_worm_x[13673:13668] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13673:13668] * PIXEL_SIZE && v_count < i_worm_y[13673:13668] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2279 < i_size && h_count >= i_worm_x[13679:13674] * PIXEL_SIZE && h_count < i_worm_x[13679:13674] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13679:13674] * PIXEL_SIZE && v_count < i_worm_y[13679:13674] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2280 < i_size && h_count >= i_worm_x[13685:13680] * PIXEL_SIZE && h_count < i_worm_x[13685:13680] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13685:13680] * PIXEL_SIZE && v_count < i_worm_y[13685:13680] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2281 < i_size && h_count >= i_worm_x[13691:13686] * PIXEL_SIZE && h_count < i_worm_x[13691:13686] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13691:13686] * PIXEL_SIZE && v_count < i_worm_y[13691:13686] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2282 < i_size && h_count >= i_worm_x[13697:13692] * PIXEL_SIZE && h_count < i_worm_x[13697:13692] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13697:13692] * PIXEL_SIZE && v_count < i_worm_y[13697:13692] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2283 < i_size && h_count >= i_worm_x[13703:13698] * PIXEL_SIZE && h_count < i_worm_x[13703:13698] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13703:13698] * PIXEL_SIZE && v_count < i_worm_y[13703:13698] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2284 < i_size && h_count >= i_worm_x[13709:13704] * PIXEL_SIZE && h_count < i_worm_x[13709:13704] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13709:13704] * PIXEL_SIZE && v_count < i_worm_y[13709:13704] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2285 < i_size && h_count >= i_worm_x[13715:13710] * PIXEL_SIZE && h_count < i_worm_x[13715:13710] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13715:13710] * PIXEL_SIZE && v_count < i_worm_y[13715:13710] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2286 < i_size && h_count >= i_worm_x[13721:13716] * PIXEL_SIZE && h_count < i_worm_x[13721:13716] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13721:13716] * PIXEL_SIZE && v_count < i_worm_y[13721:13716] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2287 < i_size && h_count >= i_worm_x[13727:13722] * PIXEL_SIZE && h_count < i_worm_x[13727:13722] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13727:13722] * PIXEL_SIZE && v_count < i_worm_y[13727:13722] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2288 < i_size && h_count >= i_worm_x[13733:13728] * PIXEL_SIZE && h_count < i_worm_x[13733:13728] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13733:13728] * PIXEL_SIZE && v_count < i_worm_y[13733:13728] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2289 < i_size && h_count >= i_worm_x[13739:13734] * PIXEL_SIZE && h_count < i_worm_x[13739:13734] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13739:13734] * PIXEL_SIZE && v_count < i_worm_y[13739:13734] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2290 < i_size && h_count >= i_worm_x[13745:13740] * PIXEL_SIZE && h_count < i_worm_x[13745:13740] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13745:13740] * PIXEL_SIZE && v_count < i_worm_y[13745:13740] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2291 < i_size && h_count >= i_worm_x[13751:13746] * PIXEL_SIZE && h_count < i_worm_x[13751:13746] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13751:13746] * PIXEL_SIZE && v_count < i_worm_y[13751:13746] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2292 < i_size && h_count >= i_worm_x[13757:13752] * PIXEL_SIZE && h_count < i_worm_x[13757:13752] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13757:13752] * PIXEL_SIZE && v_count < i_worm_y[13757:13752] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2293 < i_size && h_count >= i_worm_x[13763:13758] * PIXEL_SIZE && h_count < i_worm_x[13763:13758] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13763:13758] * PIXEL_SIZE && v_count < i_worm_y[13763:13758] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2294 < i_size && h_count >= i_worm_x[13769:13764] * PIXEL_SIZE && h_count < i_worm_x[13769:13764] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13769:13764] * PIXEL_SIZE && v_count < i_worm_y[13769:13764] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2295 < i_size && h_count >= i_worm_x[13775:13770] * PIXEL_SIZE && h_count < i_worm_x[13775:13770] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13775:13770] * PIXEL_SIZE && v_count < i_worm_y[13775:13770] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2296 < i_size && h_count >= i_worm_x[13781:13776] * PIXEL_SIZE && h_count < i_worm_x[13781:13776] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13781:13776] * PIXEL_SIZE && v_count < i_worm_y[13781:13776] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2297 < i_size && h_count >= i_worm_x[13787:13782] * PIXEL_SIZE && h_count < i_worm_x[13787:13782] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13787:13782] * PIXEL_SIZE && v_count < i_worm_y[13787:13782] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2298 < i_size && h_count >= i_worm_x[13793:13788] * PIXEL_SIZE && h_count < i_worm_x[13793:13788] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13793:13788] * PIXEL_SIZE && v_count < i_worm_y[13793:13788] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2299 < i_size && h_count >= i_worm_x[13799:13794] * PIXEL_SIZE && h_count < i_worm_x[13799:13794] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13799:13794] * PIXEL_SIZE && v_count < i_worm_y[13799:13794] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2300 < i_size && h_count >= i_worm_x[13805:13800] * PIXEL_SIZE && h_count < i_worm_x[13805:13800] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13805:13800] * PIXEL_SIZE && v_count < i_worm_y[13805:13800] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2301 < i_size && h_count >= i_worm_x[13811:13806] * PIXEL_SIZE && h_count < i_worm_x[13811:13806] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13811:13806] * PIXEL_SIZE && v_count < i_worm_y[13811:13806] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2302 < i_size && h_count >= i_worm_x[13817:13812] * PIXEL_SIZE && h_count < i_worm_x[13817:13812] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13817:13812] * PIXEL_SIZE && v_count < i_worm_y[13817:13812] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2303 < i_size && h_count >= i_worm_x[13823:13818] * PIXEL_SIZE && h_count < i_worm_x[13823:13818] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13823:13818] * PIXEL_SIZE && v_count < i_worm_y[13823:13818] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2304 < i_size && h_count >= i_worm_x[13829:13824] * PIXEL_SIZE && h_count < i_worm_x[13829:13824] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13829:13824] * PIXEL_SIZE && v_count < i_worm_y[13829:13824] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2305 < i_size && h_count >= i_worm_x[13835:13830] * PIXEL_SIZE && h_count < i_worm_x[13835:13830] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13835:13830] * PIXEL_SIZE && v_count < i_worm_y[13835:13830] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2306 < i_size && h_count >= i_worm_x[13841:13836] * PIXEL_SIZE && h_count < i_worm_x[13841:13836] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13841:13836] * PIXEL_SIZE && v_count < i_worm_y[13841:13836] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2307 < i_size && h_count >= i_worm_x[13847:13842] * PIXEL_SIZE && h_count < i_worm_x[13847:13842] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13847:13842] * PIXEL_SIZE && v_count < i_worm_y[13847:13842] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2308 < i_size && h_count >= i_worm_x[13853:13848] * PIXEL_SIZE && h_count < i_worm_x[13853:13848] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13853:13848] * PIXEL_SIZE && v_count < i_worm_y[13853:13848] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2309 < i_size && h_count >= i_worm_x[13859:13854] * PIXEL_SIZE && h_count < i_worm_x[13859:13854] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13859:13854] * PIXEL_SIZE && v_count < i_worm_y[13859:13854] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2310 < i_size && h_count >= i_worm_x[13865:13860] * PIXEL_SIZE && h_count < i_worm_x[13865:13860] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13865:13860] * PIXEL_SIZE && v_count < i_worm_y[13865:13860] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2311 < i_size && h_count >= i_worm_x[13871:13866] * PIXEL_SIZE && h_count < i_worm_x[13871:13866] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13871:13866] * PIXEL_SIZE && v_count < i_worm_y[13871:13866] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2312 < i_size && h_count >= i_worm_x[13877:13872] * PIXEL_SIZE && h_count < i_worm_x[13877:13872] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13877:13872] * PIXEL_SIZE && v_count < i_worm_y[13877:13872] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2313 < i_size && h_count >= i_worm_x[13883:13878] * PIXEL_SIZE && h_count < i_worm_x[13883:13878] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13883:13878] * PIXEL_SIZE && v_count < i_worm_y[13883:13878] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2314 < i_size && h_count >= i_worm_x[13889:13884] * PIXEL_SIZE && h_count < i_worm_x[13889:13884] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13889:13884] * PIXEL_SIZE && v_count < i_worm_y[13889:13884] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2315 < i_size && h_count >= i_worm_x[13895:13890] * PIXEL_SIZE && h_count < i_worm_x[13895:13890] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13895:13890] * PIXEL_SIZE && v_count < i_worm_y[13895:13890] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2316 < i_size && h_count >= i_worm_x[13901:13896] * PIXEL_SIZE && h_count < i_worm_x[13901:13896] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13901:13896] * PIXEL_SIZE && v_count < i_worm_y[13901:13896] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2317 < i_size && h_count >= i_worm_x[13907:13902] * PIXEL_SIZE && h_count < i_worm_x[13907:13902] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13907:13902] * PIXEL_SIZE && v_count < i_worm_y[13907:13902] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2318 < i_size && h_count >= i_worm_x[13913:13908] * PIXEL_SIZE && h_count < i_worm_x[13913:13908] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13913:13908] * PIXEL_SIZE && v_count < i_worm_y[13913:13908] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2319 < i_size && h_count >= i_worm_x[13919:13914] * PIXEL_SIZE && h_count < i_worm_x[13919:13914] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13919:13914] * PIXEL_SIZE && v_count < i_worm_y[13919:13914] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2320 < i_size && h_count >= i_worm_x[13925:13920] * PIXEL_SIZE && h_count < i_worm_x[13925:13920] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13925:13920] * PIXEL_SIZE && v_count < i_worm_y[13925:13920] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2321 < i_size && h_count >= i_worm_x[13931:13926] * PIXEL_SIZE && h_count < i_worm_x[13931:13926] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13931:13926] * PIXEL_SIZE && v_count < i_worm_y[13931:13926] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2322 < i_size && h_count >= i_worm_x[13937:13932] * PIXEL_SIZE && h_count < i_worm_x[13937:13932] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13937:13932] * PIXEL_SIZE && v_count < i_worm_y[13937:13932] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2323 < i_size && h_count >= i_worm_x[13943:13938] * PIXEL_SIZE && h_count < i_worm_x[13943:13938] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13943:13938] * PIXEL_SIZE && v_count < i_worm_y[13943:13938] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2324 < i_size && h_count >= i_worm_x[13949:13944] * PIXEL_SIZE && h_count < i_worm_x[13949:13944] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13949:13944] * PIXEL_SIZE && v_count < i_worm_y[13949:13944] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2325 < i_size && h_count >= i_worm_x[13955:13950] * PIXEL_SIZE && h_count < i_worm_x[13955:13950] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13955:13950] * PIXEL_SIZE && v_count < i_worm_y[13955:13950] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2326 < i_size && h_count >= i_worm_x[13961:13956] * PIXEL_SIZE && h_count < i_worm_x[13961:13956] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13961:13956] * PIXEL_SIZE && v_count < i_worm_y[13961:13956] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2327 < i_size && h_count >= i_worm_x[13967:13962] * PIXEL_SIZE && h_count < i_worm_x[13967:13962] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13967:13962] * PIXEL_SIZE && v_count < i_worm_y[13967:13962] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2328 < i_size && h_count >= i_worm_x[13973:13968] * PIXEL_SIZE && h_count < i_worm_x[13973:13968] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13973:13968] * PIXEL_SIZE && v_count < i_worm_y[13973:13968] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2329 < i_size && h_count >= i_worm_x[13979:13974] * PIXEL_SIZE && h_count < i_worm_x[13979:13974] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13979:13974] * PIXEL_SIZE && v_count < i_worm_y[13979:13974] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2330 < i_size && h_count >= i_worm_x[13985:13980] * PIXEL_SIZE && h_count < i_worm_x[13985:13980] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13985:13980] * PIXEL_SIZE && v_count < i_worm_y[13985:13980] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2331 < i_size && h_count >= i_worm_x[13991:13986] * PIXEL_SIZE && h_count < i_worm_x[13991:13986] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13991:13986] * PIXEL_SIZE && v_count < i_worm_y[13991:13986] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2332 < i_size && h_count >= i_worm_x[13997:13992] * PIXEL_SIZE && h_count < i_worm_x[13997:13992] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[13997:13992] * PIXEL_SIZE && v_count < i_worm_y[13997:13992] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2333 < i_size && h_count >= i_worm_x[14003:13998] * PIXEL_SIZE && h_count < i_worm_x[14003:13998] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14003:13998] * PIXEL_SIZE && v_count < i_worm_y[14003:13998] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2334 < i_size && h_count >= i_worm_x[14009:14004] * PIXEL_SIZE && h_count < i_worm_x[14009:14004] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14009:14004] * PIXEL_SIZE && v_count < i_worm_y[14009:14004] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2335 < i_size && h_count >= i_worm_x[14015:14010] * PIXEL_SIZE && h_count < i_worm_x[14015:14010] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14015:14010] * PIXEL_SIZE && v_count < i_worm_y[14015:14010] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2336 < i_size && h_count >= i_worm_x[14021:14016] * PIXEL_SIZE && h_count < i_worm_x[14021:14016] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14021:14016] * PIXEL_SIZE && v_count < i_worm_y[14021:14016] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2337 < i_size && h_count >= i_worm_x[14027:14022] * PIXEL_SIZE && h_count < i_worm_x[14027:14022] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14027:14022] * PIXEL_SIZE && v_count < i_worm_y[14027:14022] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2338 < i_size && h_count >= i_worm_x[14033:14028] * PIXEL_SIZE && h_count < i_worm_x[14033:14028] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14033:14028] * PIXEL_SIZE && v_count < i_worm_y[14033:14028] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2339 < i_size && h_count >= i_worm_x[14039:14034] * PIXEL_SIZE && h_count < i_worm_x[14039:14034] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14039:14034] * PIXEL_SIZE && v_count < i_worm_y[14039:14034] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2340 < i_size && h_count >= i_worm_x[14045:14040] * PIXEL_SIZE && h_count < i_worm_x[14045:14040] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14045:14040] * PIXEL_SIZE && v_count < i_worm_y[14045:14040] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2341 < i_size && h_count >= i_worm_x[14051:14046] * PIXEL_SIZE && h_count < i_worm_x[14051:14046] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14051:14046] * PIXEL_SIZE && v_count < i_worm_y[14051:14046] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2342 < i_size && h_count >= i_worm_x[14057:14052] * PIXEL_SIZE && h_count < i_worm_x[14057:14052] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14057:14052] * PIXEL_SIZE && v_count < i_worm_y[14057:14052] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2343 < i_size && h_count >= i_worm_x[14063:14058] * PIXEL_SIZE && h_count < i_worm_x[14063:14058] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14063:14058] * PIXEL_SIZE && v_count < i_worm_y[14063:14058] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2344 < i_size && h_count >= i_worm_x[14069:14064] * PIXEL_SIZE && h_count < i_worm_x[14069:14064] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14069:14064] * PIXEL_SIZE && v_count < i_worm_y[14069:14064] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2345 < i_size && h_count >= i_worm_x[14075:14070] * PIXEL_SIZE && h_count < i_worm_x[14075:14070] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14075:14070] * PIXEL_SIZE && v_count < i_worm_y[14075:14070] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2346 < i_size && h_count >= i_worm_x[14081:14076] * PIXEL_SIZE && h_count < i_worm_x[14081:14076] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14081:14076] * PIXEL_SIZE && v_count < i_worm_y[14081:14076] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2347 < i_size && h_count >= i_worm_x[14087:14082] * PIXEL_SIZE && h_count < i_worm_x[14087:14082] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14087:14082] * PIXEL_SIZE && v_count < i_worm_y[14087:14082] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2348 < i_size && h_count >= i_worm_x[14093:14088] * PIXEL_SIZE && h_count < i_worm_x[14093:14088] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14093:14088] * PIXEL_SIZE && v_count < i_worm_y[14093:14088] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2349 < i_size && h_count >= i_worm_x[14099:14094] * PIXEL_SIZE && h_count < i_worm_x[14099:14094] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14099:14094] * PIXEL_SIZE && v_count < i_worm_y[14099:14094] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2350 < i_size && h_count >= i_worm_x[14105:14100] * PIXEL_SIZE && h_count < i_worm_x[14105:14100] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14105:14100] * PIXEL_SIZE && v_count < i_worm_y[14105:14100] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2351 < i_size && h_count >= i_worm_x[14111:14106] * PIXEL_SIZE && h_count < i_worm_x[14111:14106] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14111:14106] * PIXEL_SIZE && v_count < i_worm_y[14111:14106] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2352 < i_size && h_count >= i_worm_x[14117:14112] * PIXEL_SIZE && h_count < i_worm_x[14117:14112] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14117:14112] * PIXEL_SIZE && v_count < i_worm_y[14117:14112] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2353 < i_size && h_count >= i_worm_x[14123:14118] * PIXEL_SIZE && h_count < i_worm_x[14123:14118] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14123:14118] * PIXEL_SIZE && v_count < i_worm_y[14123:14118] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2354 < i_size && h_count >= i_worm_x[14129:14124] * PIXEL_SIZE && h_count < i_worm_x[14129:14124] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14129:14124] * PIXEL_SIZE && v_count < i_worm_y[14129:14124] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2355 < i_size && h_count >= i_worm_x[14135:14130] * PIXEL_SIZE && h_count < i_worm_x[14135:14130] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14135:14130] * PIXEL_SIZE && v_count < i_worm_y[14135:14130] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2356 < i_size && h_count >= i_worm_x[14141:14136] * PIXEL_SIZE && h_count < i_worm_x[14141:14136] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14141:14136] * PIXEL_SIZE && v_count < i_worm_y[14141:14136] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2357 < i_size && h_count >= i_worm_x[14147:14142] * PIXEL_SIZE && h_count < i_worm_x[14147:14142] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14147:14142] * PIXEL_SIZE && v_count < i_worm_y[14147:14142] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2358 < i_size && h_count >= i_worm_x[14153:14148] * PIXEL_SIZE && h_count < i_worm_x[14153:14148] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14153:14148] * PIXEL_SIZE && v_count < i_worm_y[14153:14148] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2359 < i_size && h_count >= i_worm_x[14159:14154] * PIXEL_SIZE && h_count < i_worm_x[14159:14154] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14159:14154] * PIXEL_SIZE && v_count < i_worm_y[14159:14154] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2360 < i_size && h_count >= i_worm_x[14165:14160] * PIXEL_SIZE && h_count < i_worm_x[14165:14160] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14165:14160] * PIXEL_SIZE && v_count < i_worm_y[14165:14160] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2361 < i_size && h_count >= i_worm_x[14171:14166] * PIXEL_SIZE && h_count < i_worm_x[14171:14166] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14171:14166] * PIXEL_SIZE && v_count < i_worm_y[14171:14166] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2362 < i_size && h_count >= i_worm_x[14177:14172] * PIXEL_SIZE && h_count < i_worm_x[14177:14172] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14177:14172] * PIXEL_SIZE && v_count < i_worm_y[14177:14172] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2363 < i_size && h_count >= i_worm_x[14183:14178] * PIXEL_SIZE && h_count < i_worm_x[14183:14178] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14183:14178] * PIXEL_SIZE && v_count < i_worm_y[14183:14178] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2364 < i_size && h_count >= i_worm_x[14189:14184] * PIXEL_SIZE && h_count < i_worm_x[14189:14184] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14189:14184] * PIXEL_SIZE && v_count < i_worm_y[14189:14184] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2365 < i_size && h_count >= i_worm_x[14195:14190] * PIXEL_SIZE && h_count < i_worm_x[14195:14190] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14195:14190] * PIXEL_SIZE && v_count < i_worm_y[14195:14190] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2366 < i_size && h_count >= i_worm_x[14201:14196] * PIXEL_SIZE && h_count < i_worm_x[14201:14196] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14201:14196] * PIXEL_SIZE && v_count < i_worm_y[14201:14196] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2367 < i_size && h_count >= i_worm_x[14207:14202] * PIXEL_SIZE && h_count < i_worm_x[14207:14202] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14207:14202] * PIXEL_SIZE && v_count < i_worm_y[14207:14202] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2368 < i_size && h_count >= i_worm_x[14213:14208] * PIXEL_SIZE && h_count < i_worm_x[14213:14208] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14213:14208] * PIXEL_SIZE && v_count < i_worm_y[14213:14208] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2369 < i_size && h_count >= i_worm_x[14219:14214] * PIXEL_SIZE && h_count < i_worm_x[14219:14214] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14219:14214] * PIXEL_SIZE && v_count < i_worm_y[14219:14214] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2370 < i_size && h_count >= i_worm_x[14225:14220] * PIXEL_SIZE && h_count < i_worm_x[14225:14220] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14225:14220] * PIXEL_SIZE && v_count < i_worm_y[14225:14220] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2371 < i_size && h_count >= i_worm_x[14231:14226] * PIXEL_SIZE && h_count < i_worm_x[14231:14226] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14231:14226] * PIXEL_SIZE && v_count < i_worm_y[14231:14226] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2372 < i_size && h_count >= i_worm_x[14237:14232] * PIXEL_SIZE && h_count < i_worm_x[14237:14232] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14237:14232] * PIXEL_SIZE && v_count < i_worm_y[14237:14232] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2373 < i_size && h_count >= i_worm_x[14243:14238] * PIXEL_SIZE && h_count < i_worm_x[14243:14238] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14243:14238] * PIXEL_SIZE && v_count < i_worm_y[14243:14238] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2374 < i_size && h_count >= i_worm_x[14249:14244] * PIXEL_SIZE && h_count < i_worm_x[14249:14244] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14249:14244] * PIXEL_SIZE && v_count < i_worm_y[14249:14244] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2375 < i_size && h_count >= i_worm_x[14255:14250] * PIXEL_SIZE && h_count < i_worm_x[14255:14250] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14255:14250] * PIXEL_SIZE && v_count < i_worm_y[14255:14250] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2376 < i_size && h_count >= i_worm_x[14261:14256] * PIXEL_SIZE && h_count < i_worm_x[14261:14256] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14261:14256] * PIXEL_SIZE && v_count < i_worm_y[14261:14256] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2377 < i_size && h_count >= i_worm_x[14267:14262] * PIXEL_SIZE && h_count < i_worm_x[14267:14262] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14267:14262] * PIXEL_SIZE && v_count < i_worm_y[14267:14262] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2378 < i_size && h_count >= i_worm_x[14273:14268] * PIXEL_SIZE && h_count < i_worm_x[14273:14268] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14273:14268] * PIXEL_SIZE && v_count < i_worm_y[14273:14268] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2379 < i_size && h_count >= i_worm_x[14279:14274] * PIXEL_SIZE && h_count < i_worm_x[14279:14274] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14279:14274] * PIXEL_SIZE && v_count < i_worm_y[14279:14274] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2380 < i_size && h_count >= i_worm_x[14285:14280] * PIXEL_SIZE && h_count < i_worm_x[14285:14280] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14285:14280] * PIXEL_SIZE && v_count < i_worm_y[14285:14280] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2381 < i_size && h_count >= i_worm_x[14291:14286] * PIXEL_SIZE && h_count < i_worm_x[14291:14286] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14291:14286] * PIXEL_SIZE && v_count < i_worm_y[14291:14286] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2382 < i_size && h_count >= i_worm_x[14297:14292] * PIXEL_SIZE && h_count < i_worm_x[14297:14292] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14297:14292] * PIXEL_SIZE && v_count < i_worm_y[14297:14292] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2383 < i_size && h_count >= i_worm_x[14303:14298] * PIXEL_SIZE && h_count < i_worm_x[14303:14298] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14303:14298] * PIXEL_SIZE && v_count < i_worm_y[14303:14298] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2384 < i_size && h_count >= i_worm_x[14309:14304] * PIXEL_SIZE && h_count < i_worm_x[14309:14304] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14309:14304] * PIXEL_SIZE && v_count < i_worm_y[14309:14304] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2385 < i_size && h_count >= i_worm_x[14315:14310] * PIXEL_SIZE && h_count < i_worm_x[14315:14310] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14315:14310] * PIXEL_SIZE && v_count < i_worm_y[14315:14310] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2386 < i_size && h_count >= i_worm_x[14321:14316] * PIXEL_SIZE && h_count < i_worm_x[14321:14316] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14321:14316] * PIXEL_SIZE && v_count < i_worm_y[14321:14316] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2387 < i_size && h_count >= i_worm_x[14327:14322] * PIXEL_SIZE && h_count < i_worm_x[14327:14322] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14327:14322] * PIXEL_SIZE && v_count < i_worm_y[14327:14322] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2388 < i_size && h_count >= i_worm_x[14333:14328] * PIXEL_SIZE && h_count < i_worm_x[14333:14328] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14333:14328] * PIXEL_SIZE && v_count < i_worm_y[14333:14328] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2389 < i_size && h_count >= i_worm_x[14339:14334] * PIXEL_SIZE && h_count < i_worm_x[14339:14334] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14339:14334] * PIXEL_SIZE && v_count < i_worm_y[14339:14334] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2390 < i_size && h_count >= i_worm_x[14345:14340] * PIXEL_SIZE && h_count < i_worm_x[14345:14340] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14345:14340] * PIXEL_SIZE && v_count < i_worm_y[14345:14340] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2391 < i_size && h_count >= i_worm_x[14351:14346] * PIXEL_SIZE && h_count < i_worm_x[14351:14346] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14351:14346] * PIXEL_SIZE && v_count < i_worm_y[14351:14346] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2392 < i_size && h_count >= i_worm_x[14357:14352] * PIXEL_SIZE && h_count < i_worm_x[14357:14352] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14357:14352] * PIXEL_SIZE && v_count < i_worm_y[14357:14352] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2393 < i_size && h_count >= i_worm_x[14363:14358] * PIXEL_SIZE && h_count < i_worm_x[14363:14358] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14363:14358] * PIXEL_SIZE && v_count < i_worm_y[14363:14358] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2394 < i_size && h_count >= i_worm_x[14369:14364] * PIXEL_SIZE && h_count < i_worm_x[14369:14364] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14369:14364] * PIXEL_SIZE && v_count < i_worm_y[14369:14364] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2395 < i_size && h_count >= i_worm_x[14375:14370] * PIXEL_SIZE && h_count < i_worm_x[14375:14370] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14375:14370] * PIXEL_SIZE && v_count < i_worm_y[14375:14370] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2396 < i_size && h_count >= i_worm_x[14381:14376] * PIXEL_SIZE && h_count < i_worm_x[14381:14376] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14381:14376] * PIXEL_SIZE && v_count < i_worm_y[14381:14376] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2397 < i_size && h_count >= i_worm_x[14387:14382] * PIXEL_SIZE && h_count < i_worm_x[14387:14382] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14387:14382] * PIXEL_SIZE && v_count < i_worm_y[14387:14382] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2398 < i_size && h_count >= i_worm_x[14393:14388] * PIXEL_SIZE && h_count < i_worm_x[14393:14388] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14393:14388] * PIXEL_SIZE && v_count < i_worm_y[14393:14388] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2399 < i_size && h_count >= i_worm_x[14399:14394] * PIXEL_SIZE && h_count < i_worm_x[14399:14394] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14399:14394] * PIXEL_SIZE && v_count < i_worm_y[14399:14394] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2400 < i_size && h_count >= i_worm_x[14405:14400] * PIXEL_SIZE && h_count < i_worm_x[14405:14400] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14405:14400] * PIXEL_SIZE && v_count < i_worm_y[14405:14400] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2401 < i_size && h_count >= i_worm_x[14411:14406] * PIXEL_SIZE && h_count < i_worm_x[14411:14406] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14411:14406] * PIXEL_SIZE && v_count < i_worm_y[14411:14406] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2402 < i_size && h_count >= i_worm_x[14417:14412] * PIXEL_SIZE && h_count < i_worm_x[14417:14412] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14417:14412] * PIXEL_SIZE && v_count < i_worm_y[14417:14412] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2403 < i_size && h_count >= i_worm_x[14423:14418] * PIXEL_SIZE && h_count < i_worm_x[14423:14418] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14423:14418] * PIXEL_SIZE && v_count < i_worm_y[14423:14418] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2404 < i_size && h_count >= i_worm_x[14429:14424] * PIXEL_SIZE && h_count < i_worm_x[14429:14424] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14429:14424] * PIXEL_SIZE && v_count < i_worm_y[14429:14424] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2405 < i_size && h_count >= i_worm_x[14435:14430] * PIXEL_SIZE && h_count < i_worm_x[14435:14430] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14435:14430] * PIXEL_SIZE && v_count < i_worm_y[14435:14430] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2406 < i_size && h_count >= i_worm_x[14441:14436] * PIXEL_SIZE && h_count < i_worm_x[14441:14436] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14441:14436] * PIXEL_SIZE && v_count < i_worm_y[14441:14436] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2407 < i_size && h_count >= i_worm_x[14447:14442] * PIXEL_SIZE && h_count < i_worm_x[14447:14442] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14447:14442] * PIXEL_SIZE && v_count < i_worm_y[14447:14442] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2408 < i_size && h_count >= i_worm_x[14453:14448] * PIXEL_SIZE && h_count < i_worm_x[14453:14448] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14453:14448] * PIXEL_SIZE && v_count < i_worm_y[14453:14448] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2409 < i_size && h_count >= i_worm_x[14459:14454] * PIXEL_SIZE && h_count < i_worm_x[14459:14454] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14459:14454] * PIXEL_SIZE && v_count < i_worm_y[14459:14454] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2410 < i_size && h_count >= i_worm_x[14465:14460] * PIXEL_SIZE && h_count < i_worm_x[14465:14460] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14465:14460] * PIXEL_SIZE && v_count < i_worm_y[14465:14460] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2411 < i_size && h_count >= i_worm_x[14471:14466] * PIXEL_SIZE && h_count < i_worm_x[14471:14466] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14471:14466] * PIXEL_SIZE && v_count < i_worm_y[14471:14466] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2412 < i_size && h_count >= i_worm_x[14477:14472] * PIXEL_SIZE && h_count < i_worm_x[14477:14472] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14477:14472] * PIXEL_SIZE && v_count < i_worm_y[14477:14472] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2413 < i_size && h_count >= i_worm_x[14483:14478] * PIXEL_SIZE && h_count < i_worm_x[14483:14478] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14483:14478] * PIXEL_SIZE && v_count < i_worm_y[14483:14478] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2414 < i_size && h_count >= i_worm_x[14489:14484] * PIXEL_SIZE && h_count < i_worm_x[14489:14484] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14489:14484] * PIXEL_SIZE && v_count < i_worm_y[14489:14484] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2415 < i_size && h_count >= i_worm_x[14495:14490] * PIXEL_SIZE && h_count < i_worm_x[14495:14490] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14495:14490] * PIXEL_SIZE && v_count < i_worm_y[14495:14490] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2416 < i_size && h_count >= i_worm_x[14501:14496] * PIXEL_SIZE && h_count < i_worm_x[14501:14496] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14501:14496] * PIXEL_SIZE && v_count < i_worm_y[14501:14496] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2417 < i_size && h_count >= i_worm_x[14507:14502] * PIXEL_SIZE && h_count < i_worm_x[14507:14502] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14507:14502] * PIXEL_SIZE && v_count < i_worm_y[14507:14502] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2418 < i_size && h_count >= i_worm_x[14513:14508] * PIXEL_SIZE && h_count < i_worm_x[14513:14508] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14513:14508] * PIXEL_SIZE && v_count < i_worm_y[14513:14508] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2419 < i_size && h_count >= i_worm_x[14519:14514] * PIXEL_SIZE && h_count < i_worm_x[14519:14514] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14519:14514] * PIXEL_SIZE && v_count < i_worm_y[14519:14514] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2420 < i_size && h_count >= i_worm_x[14525:14520] * PIXEL_SIZE && h_count < i_worm_x[14525:14520] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14525:14520] * PIXEL_SIZE && v_count < i_worm_y[14525:14520] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2421 < i_size && h_count >= i_worm_x[14531:14526] * PIXEL_SIZE && h_count < i_worm_x[14531:14526] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14531:14526] * PIXEL_SIZE && v_count < i_worm_y[14531:14526] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2422 < i_size && h_count >= i_worm_x[14537:14532] * PIXEL_SIZE && h_count < i_worm_x[14537:14532] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14537:14532] * PIXEL_SIZE && v_count < i_worm_y[14537:14532] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2423 < i_size && h_count >= i_worm_x[14543:14538] * PIXEL_SIZE && h_count < i_worm_x[14543:14538] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14543:14538] * PIXEL_SIZE && v_count < i_worm_y[14543:14538] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2424 < i_size && h_count >= i_worm_x[14549:14544] * PIXEL_SIZE && h_count < i_worm_x[14549:14544] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14549:14544] * PIXEL_SIZE && v_count < i_worm_y[14549:14544] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2425 < i_size && h_count >= i_worm_x[14555:14550] * PIXEL_SIZE && h_count < i_worm_x[14555:14550] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14555:14550] * PIXEL_SIZE && v_count < i_worm_y[14555:14550] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2426 < i_size && h_count >= i_worm_x[14561:14556] * PIXEL_SIZE && h_count < i_worm_x[14561:14556] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14561:14556] * PIXEL_SIZE && v_count < i_worm_y[14561:14556] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2427 < i_size && h_count >= i_worm_x[14567:14562] * PIXEL_SIZE && h_count < i_worm_x[14567:14562] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14567:14562] * PIXEL_SIZE && v_count < i_worm_y[14567:14562] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2428 < i_size && h_count >= i_worm_x[14573:14568] * PIXEL_SIZE && h_count < i_worm_x[14573:14568] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14573:14568] * PIXEL_SIZE && v_count < i_worm_y[14573:14568] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2429 < i_size && h_count >= i_worm_x[14579:14574] * PIXEL_SIZE && h_count < i_worm_x[14579:14574] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14579:14574] * PIXEL_SIZE && v_count < i_worm_y[14579:14574] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2430 < i_size && h_count >= i_worm_x[14585:14580] * PIXEL_SIZE && h_count < i_worm_x[14585:14580] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14585:14580] * PIXEL_SIZE && v_count < i_worm_y[14585:14580] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2431 < i_size && h_count >= i_worm_x[14591:14586] * PIXEL_SIZE && h_count < i_worm_x[14591:14586] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14591:14586] * PIXEL_SIZE && v_count < i_worm_y[14591:14586] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2432 < i_size && h_count >= i_worm_x[14597:14592] * PIXEL_SIZE && h_count < i_worm_x[14597:14592] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14597:14592] * PIXEL_SIZE && v_count < i_worm_y[14597:14592] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2433 < i_size && h_count >= i_worm_x[14603:14598] * PIXEL_SIZE && h_count < i_worm_x[14603:14598] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14603:14598] * PIXEL_SIZE && v_count < i_worm_y[14603:14598] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2434 < i_size && h_count >= i_worm_x[14609:14604] * PIXEL_SIZE && h_count < i_worm_x[14609:14604] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14609:14604] * PIXEL_SIZE && v_count < i_worm_y[14609:14604] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2435 < i_size && h_count >= i_worm_x[14615:14610] * PIXEL_SIZE && h_count < i_worm_x[14615:14610] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14615:14610] * PIXEL_SIZE && v_count < i_worm_y[14615:14610] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2436 < i_size && h_count >= i_worm_x[14621:14616] * PIXEL_SIZE && h_count < i_worm_x[14621:14616] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14621:14616] * PIXEL_SIZE && v_count < i_worm_y[14621:14616] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2437 < i_size && h_count >= i_worm_x[14627:14622] * PIXEL_SIZE && h_count < i_worm_x[14627:14622] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14627:14622] * PIXEL_SIZE && v_count < i_worm_y[14627:14622] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2438 < i_size && h_count >= i_worm_x[14633:14628] * PIXEL_SIZE && h_count < i_worm_x[14633:14628] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14633:14628] * PIXEL_SIZE && v_count < i_worm_y[14633:14628] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2439 < i_size && h_count >= i_worm_x[14639:14634] * PIXEL_SIZE && h_count < i_worm_x[14639:14634] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14639:14634] * PIXEL_SIZE && v_count < i_worm_y[14639:14634] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2440 < i_size && h_count >= i_worm_x[14645:14640] * PIXEL_SIZE && h_count < i_worm_x[14645:14640] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14645:14640] * PIXEL_SIZE && v_count < i_worm_y[14645:14640] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2441 < i_size && h_count >= i_worm_x[14651:14646] * PIXEL_SIZE && h_count < i_worm_x[14651:14646] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14651:14646] * PIXEL_SIZE && v_count < i_worm_y[14651:14646] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2442 < i_size && h_count >= i_worm_x[14657:14652] * PIXEL_SIZE && h_count < i_worm_x[14657:14652] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14657:14652] * PIXEL_SIZE && v_count < i_worm_y[14657:14652] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2443 < i_size && h_count >= i_worm_x[14663:14658] * PIXEL_SIZE && h_count < i_worm_x[14663:14658] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14663:14658] * PIXEL_SIZE && v_count < i_worm_y[14663:14658] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2444 < i_size && h_count >= i_worm_x[14669:14664] * PIXEL_SIZE && h_count < i_worm_x[14669:14664] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14669:14664] * PIXEL_SIZE && v_count < i_worm_y[14669:14664] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2445 < i_size && h_count >= i_worm_x[14675:14670] * PIXEL_SIZE && h_count < i_worm_x[14675:14670] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14675:14670] * PIXEL_SIZE && v_count < i_worm_y[14675:14670] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2446 < i_size && h_count >= i_worm_x[14681:14676] * PIXEL_SIZE && h_count < i_worm_x[14681:14676] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14681:14676] * PIXEL_SIZE && v_count < i_worm_y[14681:14676] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2447 < i_size && h_count >= i_worm_x[14687:14682] * PIXEL_SIZE && h_count < i_worm_x[14687:14682] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14687:14682] * PIXEL_SIZE && v_count < i_worm_y[14687:14682] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2448 < i_size && h_count >= i_worm_x[14693:14688] * PIXEL_SIZE && h_count < i_worm_x[14693:14688] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14693:14688] * PIXEL_SIZE && v_count < i_worm_y[14693:14688] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2449 < i_size && h_count >= i_worm_x[14699:14694] * PIXEL_SIZE && h_count < i_worm_x[14699:14694] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14699:14694] * PIXEL_SIZE && v_count < i_worm_y[14699:14694] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2450 < i_size && h_count >= i_worm_x[14705:14700] * PIXEL_SIZE && h_count < i_worm_x[14705:14700] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14705:14700] * PIXEL_SIZE && v_count < i_worm_y[14705:14700] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2451 < i_size && h_count >= i_worm_x[14711:14706] * PIXEL_SIZE && h_count < i_worm_x[14711:14706] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14711:14706] * PIXEL_SIZE && v_count < i_worm_y[14711:14706] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2452 < i_size && h_count >= i_worm_x[14717:14712] * PIXEL_SIZE && h_count < i_worm_x[14717:14712] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14717:14712] * PIXEL_SIZE && v_count < i_worm_y[14717:14712] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2453 < i_size && h_count >= i_worm_x[14723:14718] * PIXEL_SIZE && h_count < i_worm_x[14723:14718] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14723:14718] * PIXEL_SIZE && v_count < i_worm_y[14723:14718] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2454 < i_size && h_count >= i_worm_x[14729:14724] * PIXEL_SIZE && h_count < i_worm_x[14729:14724] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14729:14724] * PIXEL_SIZE && v_count < i_worm_y[14729:14724] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2455 < i_size && h_count >= i_worm_x[14735:14730] * PIXEL_SIZE && h_count < i_worm_x[14735:14730] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14735:14730] * PIXEL_SIZE && v_count < i_worm_y[14735:14730] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2456 < i_size && h_count >= i_worm_x[14741:14736] * PIXEL_SIZE && h_count < i_worm_x[14741:14736] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14741:14736] * PIXEL_SIZE && v_count < i_worm_y[14741:14736] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2457 < i_size && h_count >= i_worm_x[14747:14742] * PIXEL_SIZE && h_count < i_worm_x[14747:14742] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14747:14742] * PIXEL_SIZE && v_count < i_worm_y[14747:14742] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2458 < i_size && h_count >= i_worm_x[14753:14748] * PIXEL_SIZE && h_count < i_worm_x[14753:14748] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14753:14748] * PIXEL_SIZE && v_count < i_worm_y[14753:14748] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2459 < i_size && h_count >= i_worm_x[14759:14754] * PIXEL_SIZE && h_count < i_worm_x[14759:14754] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14759:14754] * PIXEL_SIZE && v_count < i_worm_y[14759:14754] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2460 < i_size && h_count >= i_worm_x[14765:14760] * PIXEL_SIZE && h_count < i_worm_x[14765:14760] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14765:14760] * PIXEL_SIZE && v_count < i_worm_y[14765:14760] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2461 < i_size && h_count >= i_worm_x[14771:14766] * PIXEL_SIZE && h_count < i_worm_x[14771:14766] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14771:14766] * PIXEL_SIZE && v_count < i_worm_y[14771:14766] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2462 < i_size && h_count >= i_worm_x[14777:14772] * PIXEL_SIZE && h_count < i_worm_x[14777:14772] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14777:14772] * PIXEL_SIZE && v_count < i_worm_y[14777:14772] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2463 < i_size && h_count >= i_worm_x[14783:14778] * PIXEL_SIZE && h_count < i_worm_x[14783:14778] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14783:14778] * PIXEL_SIZE && v_count < i_worm_y[14783:14778] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2464 < i_size && h_count >= i_worm_x[14789:14784] * PIXEL_SIZE && h_count < i_worm_x[14789:14784] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14789:14784] * PIXEL_SIZE && v_count < i_worm_y[14789:14784] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2465 < i_size && h_count >= i_worm_x[14795:14790] * PIXEL_SIZE && h_count < i_worm_x[14795:14790] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14795:14790] * PIXEL_SIZE && v_count < i_worm_y[14795:14790] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2466 < i_size && h_count >= i_worm_x[14801:14796] * PIXEL_SIZE && h_count < i_worm_x[14801:14796] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14801:14796] * PIXEL_SIZE && v_count < i_worm_y[14801:14796] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2467 < i_size && h_count >= i_worm_x[14807:14802] * PIXEL_SIZE && h_count < i_worm_x[14807:14802] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14807:14802] * PIXEL_SIZE && v_count < i_worm_y[14807:14802] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2468 < i_size && h_count >= i_worm_x[14813:14808] * PIXEL_SIZE && h_count < i_worm_x[14813:14808] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14813:14808] * PIXEL_SIZE && v_count < i_worm_y[14813:14808] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2469 < i_size && h_count >= i_worm_x[14819:14814] * PIXEL_SIZE && h_count < i_worm_x[14819:14814] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14819:14814] * PIXEL_SIZE && v_count < i_worm_y[14819:14814] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2470 < i_size && h_count >= i_worm_x[14825:14820] * PIXEL_SIZE && h_count < i_worm_x[14825:14820] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14825:14820] * PIXEL_SIZE && v_count < i_worm_y[14825:14820] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2471 < i_size && h_count >= i_worm_x[14831:14826] * PIXEL_SIZE && h_count < i_worm_x[14831:14826] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14831:14826] * PIXEL_SIZE && v_count < i_worm_y[14831:14826] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2472 < i_size && h_count >= i_worm_x[14837:14832] * PIXEL_SIZE && h_count < i_worm_x[14837:14832] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14837:14832] * PIXEL_SIZE && v_count < i_worm_y[14837:14832] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2473 < i_size && h_count >= i_worm_x[14843:14838] * PIXEL_SIZE && h_count < i_worm_x[14843:14838] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14843:14838] * PIXEL_SIZE && v_count < i_worm_y[14843:14838] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2474 < i_size && h_count >= i_worm_x[14849:14844] * PIXEL_SIZE && h_count < i_worm_x[14849:14844] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14849:14844] * PIXEL_SIZE && v_count < i_worm_y[14849:14844] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2475 < i_size && h_count >= i_worm_x[14855:14850] * PIXEL_SIZE && h_count < i_worm_x[14855:14850] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14855:14850] * PIXEL_SIZE && v_count < i_worm_y[14855:14850] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2476 < i_size && h_count >= i_worm_x[14861:14856] * PIXEL_SIZE && h_count < i_worm_x[14861:14856] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14861:14856] * PIXEL_SIZE && v_count < i_worm_y[14861:14856] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2477 < i_size && h_count >= i_worm_x[14867:14862] * PIXEL_SIZE && h_count < i_worm_x[14867:14862] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14867:14862] * PIXEL_SIZE && v_count < i_worm_y[14867:14862] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2478 < i_size && h_count >= i_worm_x[14873:14868] * PIXEL_SIZE && h_count < i_worm_x[14873:14868] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14873:14868] * PIXEL_SIZE && v_count < i_worm_y[14873:14868] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2479 < i_size && h_count >= i_worm_x[14879:14874] * PIXEL_SIZE && h_count < i_worm_x[14879:14874] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14879:14874] * PIXEL_SIZE && v_count < i_worm_y[14879:14874] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2480 < i_size && h_count >= i_worm_x[14885:14880] * PIXEL_SIZE && h_count < i_worm_x[14885:14880] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14885:14880] * PIXEL_SIZE && v_count < i_worm_y[14885:14880] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2481 < i_size && h_count >= i_worm_x[14891:14886] * PIXEL_SIZE && h_count < i_worm_x[14891:14886] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14891:14886] * PIXEL_SIZE && v_count < i_worm_y[14891:14886] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2482 < i_size && h_count >= i_worm_x[14897:14892] * PIXEL_SIZE && h_count < i_worm_x[14897:14892] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14897:14892] * PIXEL_SIZE && v_count < i_worm_y[14897:14892] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2483 < i_size && h_count >= i_worm_x[14903:14898] * PIXEL_SIZE && h_count < i_worm_x[14903:14898] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14903:14898] * PIXEL_SIZE && v_count < i_worm_y[14903:14898] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2484 < i_size && h_count >= i_worm_x[14909:14904] * PIXEL_SIZE && h_count < i_worm_x[14909:14904] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14909:14904] * PIXEL_SIZE && v_count < i_worm_y[14909:14904] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2485 < i_size && h_count >= i_worm_x[14915:14910] * PIXEL_SIZE && h_count < i_worm_x[14915:14910] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14915:14910] * PIXEL_SIZE && v_count < i_worm_y[14915:14910] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2486 < i_size && h_count >= i_worm_x[14921:14916] * PIXEL_SIZE && h_count < i_worm_x[14921:14916] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14921:14916] * PIXEL_SIZE && v_count < i_worm_y[14921:14916] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2487 < i_size && h_count >= i_worm_x[14927:14922] * PIXEL_SIZE && h_count < i_worm_x[14927:14922] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14927:14922] * PIXEL_SIZE && v_count < i_worm_y[14927:14922] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2488 < i_size && h_count >= i_worm_x[14933:14928] * PIXEL_SIZE && h_count < i_worm_x[14933:14928] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14933:14928] * PIXEL_SIZE && v_count < i_worm_y[14933:14928] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2489 < i_size && h_count >= i_worm_x[14939:14934] * PIXEL_SIZE && h_count < i_worm_x[14939:14934] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14939:14934] * PIXEL_SIZE && v_count < i_worm_y[14939:14934] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2490 < i_size && h_count >= i_worm_x[14945:14940] * PIXEL_SIZE && h_count < i_worm_x[14945:14940] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14945:14940] * PIXEL_SIZE && v_count < i_worm_y[14945:14940] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2491 < i_size && h_count >= i_worm_x[14951:14946] * PIXEL_SIZE && h_count < i_worm_x[14951:14946] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14951:14946] * PIXEL_SIZE && v_count < i_worm_y[14951:14946] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2492 < i_size && h_count >= i_worm_x[14957:14952] * PIXEL_SIZE && h_count < i_worm_x[14957:14952] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14957:14952] * PIXEL_SIZE && v_count < i_worm_y[14957:14952] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2493 < i_size && h_count >= i_worm_x[14963:14958] * PIXEL_SIZE && h_count < i_worm_x[14963:14958] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14963:14958] * PIXEL_SIZE && v_count < i_worm_y[14963:14958] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2494 < i_size && h_count >= i_worm_x[14969:14964] * PIXEL_SIZE && h_count < i_worm_x[14969:14964] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14969:14964] * PIXEL_SIZE && v_count < i_worm_y[14969:14964] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2495 < i_size && h_count >= i_worm_x[14975:14970] * PIXEL_SIZE && h_count < i_worm_x[14975:14970] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14975:14970] * PIXEL_SIZE && v_count < i_worm_y[14975:14970] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2496 < i_size && h_count >= i_worm_x[14981:14976] * PIXEL_SIZE && h_count < i_worm_x[14981:14976] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14981:14976] * PIXEL_SIZE && v_count < i_worm_y[14981:14976] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2497 < i_size && h_count >= i_worm_x[14987:14982] * PIXEL_SIZE && h_count < i_worm_x[14987:14982] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14987:14982] * PIXEL_SIZE && v_count < i_worm_y[14987:14982] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2498 < i_size && h_count >= i_worm_x[14993:14988] * PIXEL_SIZE && h_count < i_worm_x[14993:14988] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14993:14988] * PIXEL_SIZE && v_count < i_worm_y[14993:14988] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2499 < i_size && h_count >= i_worm_x[14999:14994] * PIXEL_SIZE && h_count < i_worm_x[14999:14994] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[14999:14994] * PIXEL_SIZE && v_count < i_worm_y[14999:14994] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2500 < i_size && h_count >= i_worm_x[15005:15000] * PIXEL_SIZE && h_count < i_worm_x[15005:15000] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15005:15000] * PIXEL_SIZE && v_count < i_worm_y[15005:15000] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2501 < i_size && h_count >= i_worm_x[15011:15006] * PIXEL_SIZE && h_count < i_worm_x[15011:15006] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15011:15006] * PIXEL_SIZE && v_count < i_worm_y[15011:15006] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2502 < i_size && h_count >= i_worm_x[15017:15012] * PIXEL_SIZE && h_count < i_worm_x[15017:15012] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15017:15012] * PIXEL_SIZE && v_count < i_worm_y[15017:15012] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2503 < i_size && h_count >= i_worm_x[15023:15018] * PIXEL_SIZE && h_count < i_worm_x[15023:15018] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15023:15018] * PIXEL_SIZE && v_count < i_worm_y[15023:15018] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2504 < i_size && h_count >= i_worm_x[15029:15024] * PIXEL_SIZE && h_count < i_worm_x[15029:15024] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15029:15024] * PIXEL_SIZE && v_count < i_worm_y[15029:15024] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2505 < i_size && h_count >= i_worm_x[15035:15030] * PIXEL_SIZE && h_count < i_worm_x[15035:15030] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15035:15030] * PIXEL_SIZE && v_count < i_worm_y[15035:15030] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2506 < i_size && h_count >= i_worm_x[15041:15036] * PIXEL_SIZE && h_count < i_worm_x[15041:15036] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15041:15036] * PIXEL_SIZE && v_count < i_worm_y[15041:15036] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2507 < i_size && h_count >= i_worm_x[15047:15042] * PIXEL_SIZE && h_count < i_worm_x[15047:15042] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15047:15042] * PIXEL_SIZE && v_count < i_worm_y[15047:15042] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2508 < i_size && h_count >= i_worm_x[15053:15048] * PIXEL_SIZE && h_count < i_worm_x[15053:15048] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15053:15048] * PIXEL_SIZE && v_count < i_worm_y[15053:15048] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2509 < i_size && h_count >= i_worm_x[15059:15054] * PIXEL_SIZE && h_count < i_worm_x[15059:15054] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15059:15054] * PIXEL_SIZE && v_count < i_worm_y[15059:15054] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2510 < i_size && h_count >= i_worm_x[15065:15060] * PIXEL_SIZE && h_count < i_worm_x[15065:15060] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15065:15060] * PIXEL_SIZE && v_count < i_worm_y[15065:15060] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2511 < i_size && h_count >= i_worm_x[15071:15066] * PIXEL_SIZE && h_count < i_worm_x[15071:15066] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15071:15066] * PIXEL_SIZE && v_count < i_worm_y[15071:15066] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2512 < i_size && h_count >= i_worm_x[15077:15072] * PIXEL_SIZE && h_count < i_worm_x[15077:15072] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15077:15072] * PIXEL_SIZE && v_count < i_worm_y[15077:15072] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2513 < i_size && h_count >= i_worm_x[15083:15078] * PIXEL_SIZE && h_count < i_worm_x[15083:15078] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15083:15078] * PIXEL_SIZE && v_count < i_worm_y[15083:15078] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2514 < i_size && h_count >= i_worm_x[15089:15084] * PIXEL_SIZE && h_count < i_worm_x[15089:15084] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15089:15084] * PIXEL_SIZE && v_count < i_worm_y[15089:15084] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2515 < i_size && h_count >= i_worm_x[15095:15090] * PIXEL_SIZE && h_count < i_worm_x[15095:15090] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15095:15090] * PIXEL_SIZE && v_count < i_worm_y[15095:15090] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2516 < i_size && h_count >= i_worm_x[15101:15096] * PIXEL_SIZE && h_count < i_worm_x[15101:15096] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15101:15096] * PIXEL_SIZE && v_count < i_worm_y[15101:15096] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2517 < i_size && h_count >= i_worm_x[15107:15102] * PIXEL_SIZE && h_count < i_worm_x[15107:15102] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15107:15102] * PIXEL_SIZE && v_count < i_worm_y[15107:15102] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2518 < i_size && h_count >= i_worm_x[15113:15108] * PIXEL_SIZE && h_count < i_worm_x[15113:15108] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15113:15108] * PIXEL_SIZE && v_count < i_worm_y[15113:15108] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2519 < i_size && h_count >= i_worm_x[15119:15114] * PIXEL_SIZE && h_count < i_worm_x[15119:15114] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15119:15114] * PIXEL_SIZE && v_count < i_worm_y[15119:15114] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2520 < i_size && h_count >= i_worm_x[15125:15120] * PIXEL_SIZE && h_count < i_worm_x[15125:15120] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15125:15120] * PIXEL_SIZE && v_count < i_worm_y[15125:15120] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2521 < i_size && h_count >= i_worm_x[15131:15126] * PIXEL_SIZE && h_count < i_worm_x[15131:15126] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15131:15126] * PIXEL_SIZE && v_count < i_worm_y[15131:15126] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2522 < i_size && h_count >= i_worm_x[15137:15132] * PIXEL_SIZE && h_count < i_worm_x[15137:15132] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15137:15132] * PIXEL_SIZE && v_count < i_worm_y[15137:15132] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2523 < i_size && h_count >= i_worm_x[15143:15138] * PIXEL_SIZE && h_count < i_worm_x[15143:15138] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15143:15138] * PIXEL_SIZE && v_count < i_worm_y[15143:15138] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2524 < i_size && h_count >= i_worm_x[15149:15144] * PIXEL_SIZE && h_count < i_worm_x[15149:15144] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15149:15144] * PIXEL_SIZE && v_count < i_worm_y[15149:15144] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2525 < i_size && h_count >= i_worm_x[15155:15150] * PIXEL_SIZE && h_count < i_worm_x[15155:15150] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15155:15150] * PIXEL_SIZE && v_count < i_worm_y[15155:15150] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2526 < i_size && h_count >= i_worm_x[15161:15156] * PIXEL_SIZE && h_count < i_worm_x[15161:15156] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15161:15156] * PIXEL_SIZE && v_count < i_worm_y[15161:15156] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2527 < i_size && h_count >= i_worm_x[15167:15162] * PIXEL_SIZE && h_count < i_worm_x[15167:15162] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15167:15162] * PIXEL_SIZE && v_count < i_worm_y[15167:15162] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2528 < i_size && h_count >= i_worm_x[15173:15168] * PIXEL_SIZE && h_count < i_worm_x[15173:15168] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15173:15168] * PIXEL_SIZE && v_count < i_worm_y[15173:15168] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2529 < i_size && h_count >= i_worm_x[15179:15174] * PIXEL_SIZE && h_count < i_worm_x[15179:15174] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15179:15174] * PIXEL_SIZE && v_count < i_worm_y[15179:15174] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2530 < i_size && h_count >= i_worm_x[15185:15180] * PIXEL_SIZE && h_count < i_worm_x[15185:15180] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15185:15180] * PIXEL_SIZE && v_count < i_worm_y[15185:15180] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2531 < i_size && h_count >= i_worm_x[15191:15186] * PIXEL_SIZE && h_count < i_worm_x[15191:15186] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15191:15186] * PIXEL_SIZE && v_count < i_worm_y[15191:15186] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2532 < i_size && h_count >= i_worm_x[15197:15192] * PIXEL_SIZE && h_count < i_worm_x[15197:15192] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15197:15192] * PIXEL_SIZE && v_count < i_worm_y[15197:15192] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2533 < i_size && h_count >= i_worm_x[15203:15198] * PIXEL_SIZE && h_count < i_worm_x[15203:15198] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15203:15198] * PIXEL_SIZE && v_count < i_worm_y[15203:15198] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2534 < i_size && h_count >= i_worm_x[15209:15204] * PIXEL_SIZE && h_count < i_worm_x[15209:15204] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15209:15204] * PIXEL_SIZE && v_count < i_worm_y[15209:15204] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2535 < i_size && h_count >= i_worm_x[15215:15210] * PIXEL_SIZE && h_count < i_worm_x[15215:15210] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15215:15210] * PIXEL_SIZE && v_count < i_worm_y[15215:15210] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2536 < i_size && h_count >= i_worm_x[15221:15216] * PIXEL_SIZE && h_count < i_worm_x[15221:15216] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15221:15216] * PIXEL_SIZE && v_count < i_worm_y[15221:15216] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2537 < i_size && h_count >= i_worm_x[15227:15222] * PIXEL_SIZE && h_count < i_worm_x[15227:15222] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15227:15222] * PIXEL_SIZE && v_count < i_worm_y[15227:15222] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2538 < i_size && h_count >= i_worm_x[15233:15228] * PIXEL_SIZE && h_count < i_worm_x[15233:15228] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15233:15228] * PIXEL_SIZE && v_count < i_worm_y[15233:15228] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2539 < i_size && h_count >= i_worm_x[15239:15234] * PIXEL_SIZE && h_count < i_worm_x[15239:15234] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15239:15234] * PIXEL_SIZE && v_count < i_worm_y[15239:15234] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2540 < i_size && h_count >= i_worm_x[15245:15240] * PIXEL_SIZE && h_count < i_worm_x[15245:15240] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15245:15240] * PIXEL_SIZE && v_count < i_worm_y[15245:15240] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2541 < i_size && h_count >= i_worm_x[15251:15246] * PIXEL_SIZE && h_count < i_worm_x[15251:15246] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15251:15246] * PIXEL_SIZE && v_count < i_worm_y[15251:15246] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2542 < i_size && h_count >= i_worm_x[15257:15252] * PIXEL_SIZE && h_count < i_worm_x[15257:15252] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15257:15252] * PIXEL_SIZE && v_count < i_worm_y[15257:15252] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2543 < i_size && h_count >= i_worm_x[15263:15258] * PIXEL_SIZE && h_count < i_worm_x[15263:15258] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15263:15258] * PIXEL_SIZE && v_count < i_worm_y[15263:15258] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2544 < i_size && h_count >= i_worm_x[15269:15264] * PIXEL_SIZE && h_count < i_worm_x[15269:15264] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15269:15264] * PIXEL_SIZE && v_count < i_worm_y[15269:15264] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2545 < i_size && h_count >= i_worm_x[15275:15270] * PIXEL_SIZE && h_count < i_worm_x[15275:15270] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15275:15270] * PIXEL_SIZE && v_count < i_worm_y[15275:15270] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2546 < i_size && h_count >= i_worm_x[15281:15276] * PIXEL_SIZE && h_count < i_worm_x[15281:15276] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15281:15276] * PIXEL_SIZE && v_count < i_worm_y[15281:15276] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2547 < i_size && h_count >= i_worm_x[15287:15282] * PIXEL_SIZE && h_count < i_worm_x[15287:15282] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15287:15282] * PIXEL_SIZE && v_count < i_worm_y[15287:15282] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2548 < i_size && h_count >= i_worm_x[15293:15288] * PIXEL_SIZE && h_count < i_worm_x[15293:15288] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15293:15288] * PIXEL_SIZE && v_count < i_worm_y[15293:15288] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2549 < i_size && h_count >= i_worm_x[15299:15294] * PIXEL_SIZE && h_count < i_worm_x[15299:15294] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15299:15294] * PIXEL_SIZE && v_count < i_worm_y[15299:15294] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2550 < i_size && h_count >= i_worm_x[15305:15300] * PIXEL_SIZE && h_count < i_worm_x[15305:15300] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15305:15300] * PIXEL_SIZE && v_count < i_worm_y[15305:15300] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2551 < i_size && h_count >= i_worm_x[15311:15306] * PIXEL_SIZE && h_count < i_worm_x[15311:15306] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15311:15306] * PIXEL_SIZE && v_count < i_worm_y[15311:15306] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2552 < i_size && h_count >= i_worm_x[15317:15312] * PIXEL_SIZE && h_count < i_worm_x[15317:15312] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15317:15312] * PIXEL_SIZE && v_count < i_worm_y[15317:15312] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2553 < i_size && h_count >= i_worm_x[15323:15318] * PIXEL_SIZE && h_count < i_worm_x[15323:15318] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15323:15318] * PIXEL_SIZE && v_count < i_worm_y[15323:15318] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2554 < i_size && h_count >= i_worm_x[15329:15324] * PIXEL_SIZE && h_count < i_worm_x[15329:15324] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15329:15324] * PIXEL_SIZE && v_count < i_worm_y[15329:15324] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2555 < i_size && h_count >= i_worm_x[15335:15330] * PIXEL_SIZE && h_count < i_worm_x[15335:15330] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15335:15330] * PIXEL_SIZE && v_count < i_worm_y[15335:15330] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2556 < i_size && h_count >= i_worm_x[15341:15336] * PIXEL_SIZE && h_count < i_worm_x[15341:15336] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15341:15336] * PIXEL_SIZE && v_count < i_worm_y[15341:15336] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2557 < i_size && h_count >= i_worm_x[15347:15342] * PIXEL_SIZE && h_count < i_worm_x[15347:15342] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15347:15342] * PIXEL_SIZE && v_count < i_worm_y[15347:15342] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2558 < i_size && h_count >= i_worm_x[15353:15348] * PIXEL_SIZE && h_count < i_worm_x[15353:15348] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15353:15348] * PIXEL_SIZE && v_count < i_worm_y[15353:15348] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2559 < i_size && h_count >= i_worm_x[15359:15354] * PIXEL_SIZE && h_count < i_worm_x[15359:15354] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15359:15354] * PIXEL_SIZE && v_count < i_worm_y[15359:15354] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2560 < i_size && h_count >= i_worm_x[15365:15360] * PIXEL_SIZE && h_count < i_worm_x[15365:15360] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15365:15360] * PIXEL_SIZE && v_count < i_worm_y[15365:15360] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2561 < i_size && h_count >= i_worm_x[15371:15366] * PIXEL_SIZE && h_count < i_worm_x[15371:15366] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15371:15366] * PIXEL_SIZE && v_count < i_worm_y[15371:15366] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2562 < i_size && h_count >= i_worm_x[15377:15372] * PIXEL_SIZE && h_count < i_worm_x[15377:15372] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15377:15372] * PIXEL_SIZE && v_count < i_worm_y[15377:15372] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2563 < i_size && h_count >= i_worm_x[15383:15378] * PIXEL_SIZE && h_count < i_worm_x[15383:15378] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15383:15378] * PIXEL_SIZE && v_count < i_worm_y[15383:15378] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2564 < i_size && h_count >= i_worm_x[15389:15384] * PIXEL_SIZE && h_count < i_worm_x[15389:15384] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15389:15384] * PIXEL_SIZE && v_count < i_worm_y[15389:15384] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2565 < i_size && h_count >= i_worm_x[15395:15390] * PIXEL_SIZE && h_count < i_worm_x[15395:15390] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15395:15390] * PIXEL_SIZE && v_count < i_worm_y[15395:15390] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2566 < i_size && h_count >= i_worm_x[15401:15396] * PIXEL_SIZE && h_count < i_worm_x[15401:15396] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15401:15396] * PIXEL_SIZE && v_count < i_worm_y[15401:15396] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2567 < i_size && h_count >= i_worm_x[15407:15402] * PIXEL_SIZE && h_count < i_worm_x[15407:15402] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15407:15402] * PIXEL_SIZE && v_count < i_worm_y[15407:15402] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2568 < i_size && h_count >= i_worm_x[15413:15408] * PIXEL_SIZE && h_count < i_worm_x[15413:15408] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15413:15408] * PIXEL_SIZE && v_count < i_worm_y[15413:15408] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2569 < i_size && h_count >= i_worm_x[15419:15414] * PIXEL_SIZE && h_count < i_worm_x[15419:15414] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15419:15414] * PIXEL_SIZE && v_count < i_worm_y[15419:15414] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2570 < i_size && h_count >= i_worm_x[15425:15420] * PIXEL_SIZE && h_count < i_worm_x[15425:15420] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15425:15420] * PIXEL_SIZE && v_count < i_worm_y[15425:15420] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2571 < i_size && h_count >= i_worm_x[15431:15426] * PIXEL_SIZE && h_count < i_worm_x[15431:15426] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15431:15426] * PIXEL_SIZE && v_count < i_worm_y[15431:15426] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2572 < i_size && h_count >= i_worm_x[15437:15432] * PIXEL_SIZE && h_count < i_worm_x[15437:15432] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15437:15432] * PIXEL_SIZE && v_count < i_worm_y[15437:15432] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2573 < i_size && h_count >= i_worm_x[15443:15438] * PIXEL_SIZE && h_count < i_worm_x[15443:15438] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15443:15438] * PIXEL_SIZE && v_count < i_worm_y[15443:15438] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2574 < i_size && h_count >= i_worm_x[15449:15444] * PIXEL_SIZE && h_count < i_worm_x[15449:15444] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15449:15444] * PIXEL_SIZE && v_count < i_worm_y[15449:15444] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2575 < i_size && h_count >= i_worm_x[15455:15450] * PIXEL_SIZE && h_count < i_worm_x[15455:15450] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15455:15450] * PIXEL_SIZE && v_count < i_worm_y[15455:15450] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2576 < i_size && h_count >= i_worm_x[15461:15456] * PIXEL_SIZE && h_count < i_worm_x[15461:15456] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15461:15456] * PIXEL_SIZE && v_count < i_worm_y[15461:15456] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2577 < i_size && h_count >= i_worm_x[15467:15462] * PIXEL_SIZE && h_count < i_worm_x[15467:15462] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15467:15462] * PIXEL_SIZE && v_count < i_worm_y[15467:15462] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2578 < i_size && h_count >= i_worm_x[15473:15468] * PIXEL_SIZE && h_count < i_worm_x[15473:15468] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15473:15468] * PIXEL_SIZE && v_count < i_worm_y[15473:15468] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2579 < i_size && h_count >= i_worm_x[15479:15474] * PIXEL_SIZE && h_count < i_worm_x[15479:15474] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15479:15474] * PIXEL_SIZE && v_count < i_worm_y[15479:15474] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2580 < i_size && h_count >= i_worm_x[15485:15480] * PIXEL_SIZE && h_count < i_worm_x[15485:15480] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15485:15480] * PIXEL_SIZE && v_count < i_worm_y[15485:15480] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2581 < i_size && h_count >= i_worm_x[15491:15486] * PIXEL_SIZE && h_count < i_worm_x[15491:15486] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15491:15486] * PIXEL_SIZE && v_count < i_worm_y[15491:15486] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2582 < i_size && h_count >= i_worm_x[15497:15492] * PIXEL_SIZE && h_count < i_worm_x[15497:15492] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15497:15492] * PIXEL_SIZE && v_count < i_worm_y[15497:15492] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2583 < i_size && h_count >= i_worm_x[15503:15498] * PIXEL_SIZE && h_count < i_worm_x[15503:15498] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15503:15498] * PIXEL_SIZE && v_count < i_worm_y[15503:15498] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2584 < i_size && h_count >= i_worm_x[15509:15504] * PIXEL_SIZE && h_count < i_worm_x[15509:15504] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15509:15504] * PIXEL_SIZE && v_count < i_worm_y[15509:15504] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2585 < i_size && h_count >= i_worm_x[15515:15510] * PIXEL_SIZE && h_count < i_worm_x[15515:15510] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15515:15510] * PIXEL_SIZE && v_count < i_worm_y[15515:15510] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2586 < i_size && h_count >= i_worm_x[15521:15516] * PIXEL_SIZE && h_count < i_worm_x[15521:15516] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15521:15516] * PIXEL_SIZE && v_count < i_worm_y[15521:15516] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2587 < i_size && h_count >= i_worm_x[15527:15522] * PIXEL_SIZE && h_count < i_worm_x[15527:15522] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15527:15522] * PIXEL_SIZE && v_count < i_worm_y[15527:15522] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2588 < i_size && h_count >= i_worm_x[15533:15528] * PIXEL_SIZE && h_count < i_worm_x[15533:15528] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15533:15528] * PIXEL_SIZE && v_count < i_worm_y[15533:15528] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2589 < i_size && h_count >= i_worm_x[15539:15534] * PIXEL_SIZE && h_count < i_worm_x[15539:15534] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15539:15534] * PIXEL_SIZE && v_count < i_worm_y[15539:15534] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2590 < i_size && h_count >= i_worm_x[15545:15540] * PIXEL_SIZE && h_count < i_worm_x[15545:15540] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15545:15540] * PIXEL_SIZE && v_count < i_worm_y[15545:15540] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2591 < i_size && h_count >= i_worm_x[15551:15546] * PIXEL_SIZE && h_count < i_worm_x[15551:15546] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15551:15546] * PIXEL_SIZE && v_count < i_worm_y[15551:15546] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2592 < i_size && h_count >= i_worm_x[15557:15552] * PIXEL_SIZE && h_count < i_worm_x[15557:15552] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15557:15552] * PIXEL_SIZE && v_count < i_worm_y[15557:15552] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2593 < i_size && h_count >= i_worm_x[15563:15558] * PIXEL_SIZE && h_count < i_worm_x[15563:15558] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15563:15558] * PIXEL_SIZE && v_count < i_worm_y[15563:15558] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2594 < i_size && h_count >= i_worm_x[15569:15564] * PIXEL_SIZE && h_count < i_worm_x[15569:15564] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15569:15564] * PIXEL_SIZE && v_count < i_worm_y[15569:15564] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2595 < i_size && h_count >= i_worm_x[15575:15570] * PIXEL_SIZE && h_count < i_worm_x[15575:15570] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15575:15570] * PIXEL_SIZE && v_count < i_worm_y[15575:15570] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2596 < i_size && h_count >= i_worm_x[15581:15576] * PIXEL_SIZE && h_count < i_worm_x[15581:15576] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15581:15576] * PIXEL_SIZE && v_count < i_worm_y[15581:15576] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2597 < i_size && h_count >= i_worm_x[15587:15582] * PIXEL_SIZE && h_count < i_worm_x[15587:15582] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15587:15582] * PIXEL_SIZE && v_count < i_worm_y[15587:15582] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2598 < i_size && h_count >= i_worm_x[15593:15588] * PIXEL_SIZE && h_count < i_worm_x[15593:15588] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15593:15588] * PIXEL_SIZE && v_count < i_worm_y[15593:15588] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2599 < i_size && h_count >= i_worm_x[15599:15594] * PIXEL_SIZE && h_count < i_worm_x[15599:15594] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15599:15594] * PIXEL_SIZE && v_count < i_worm_y[15599:15594] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2600 < i_size && h_count >= i_worm_x[15605:15600] * PIXEL_SIZE && h_count < i_worm_x[15605:15600] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15605:15600] * PIXEL_SIZE && v_count < i_worm_y[15605:15600] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2601 < i_size && h_count >= i_worm_x[15611:15606] * PIXEL_SIZE && h_count < i_worm_x[15611:15606] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15611:15606] * PIXEL_SIZE && v_count < i_worm_y[15611:15606] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2602 < i_size && h_count >= i_worm_x[15617:15612] * PIXEL_SIZE && h_count < i_worm_x[15617:15612] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15617:15612] * PIXEL_SIZE && v_count < i_worm_y[15617:15612] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2603 < i_size && h_count >= i_worm_x[15623:15618] * PIXEL_SIZE && h_count < i_worm_x[15623:15618] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15623:15618] * PIXEL_SIZE && v_count < i_worm_y[15623:15618] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2604 < i_size && h_count >= i_worm_x[15629:15624] * PIXEL_SIZE && h_count < i_worm_x[15629:15624] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15629:15624] * PIXEL_SIZE && v_count < i_worm_y[15629:15624] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2605 < i_size && h_count >= i_worm_x[15635:15630] * PIXEL_SIZE && h_count < i_worm_x[15635:15630] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15635:15630] * PIXEL_SIZE && v_count < i_worm_y[15635:15630] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2606 < i_size && h_count >= i_worm_x[15641:15636] * PIXEL_SIZE && h_count < i_worm_x[15641:15636] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15641:15636] * PIXEL_SIZE && v_count < i_worm_y[15641:15636] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2607 < i_size && h_count >= i_worm_x[15647:15642] * PIXEL_SIZE && h_count < i_worm_x[15647:15642] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15647:15642] * PIXEL_SIZE && v_count < i_worm_y[15647:15642] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2608 < i_size && h_count >= i_worm_x[15653:15648] * PIXEL_SIZE && h_count < i_worm_x[15653:15648] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15653:15648] * PIXEL_SIZE && v_count < i_worm_y[15653:15648] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2609 < i_size && h_count >= i_worm_x[15659:15654] * PIXEL_SIZE && h_count < i_worm_x[15659:15654] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15659:15654] * PIXEL_SIZE && v_count < i_worm_y[15659:15654] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2610 < i_size && h_count >= i_worm_x[15665:15660] * PIXEL_SIZE && h_count < i_worm_x[15665:15660] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15665:15660] * PIXEL_SIZE && v_count < i_worm_y[15665:15660] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2611 < i_size && h_count >= i_worm_x[15671:15666] * PIXEL_SIZE && h_count < i_worm_x[15671:15666] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15671:15666] * PIXEL_SIZE && v_count < i_worm_y[15671:15666] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2612 < i_size && h_count >= i_worm_x[15677:15672] * PIXEL_SIZE && h_count < i_worm_x[15677:15672] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15677:15672] * PIXEL_SIZE && v_count < i_worm_y[15677:15672] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2613 < i_size && h_count >= i_worm_x[15683:15678] * PIXEL_SIZE && h_count < i_worm_x[15683:15678] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15683:15678] * PIXEL_SIZE && v_count < i_worm_y[15683:15678] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2614 < i_size && h_count >= i_worm_x[15689:15684] * PIXEL_SIZE && h_count < i_worm_x[15689:15684] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15689:15684] * PIXEL_SIZE && v_count < i_worm_y[15689:15684] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2615 < i_size && h_count >= i_worm_x[15695:15690] * PIXEL_SIZE && h_count < i_worm_x[15695:15690] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15695:15690] * PIXEL_SIZE && v_count < i_worm_y[15695:15690] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2616 < i_size && h_count >= i_worm_x[15701:15696] * PIXEL_SIZE && h_count < i_worm_x[15701:15696] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15701:15696] * PIXEL_SIZE && v_count < i_worm_y[15701:15696] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2617 < i_size && h_count >= i_worm_x[15707:15702] * PIXEL_SIZE && h_count < i_worm_x[15707:15702] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15707:15702] * PIXEL_SIZE && v_count < i_worm_y[15707:15702] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2618 < i_size && h_count >= i_worm_x[15713:15708] * PIXEL_SIZE && h_count < i_worm_x[15713:15708] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15713:15708] * PIXEL_SIZE && v_count < i_worm_y[15713:15708] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2619 < i_size && h_count >= i_worm_x[15719:15714] * PIXEL_SIZE && h_count < i_worm_x[15719:15714] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15719:15714] * PIXEL_SIZE && v_count < i_worm_y[15719:15714] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2620 < i_size && h_count >= i_worm_x[15725:15720] * PIXEL_SIZE && h_count < i_worm_x[15725:15720] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15725:15720] * PIXEL_SIZE && v_count < i_worm_y[15725:15720] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2621 < i_size && h_count >= i_worm_x[15731:15726] * PIXEL_SIZE && h_count < i_worm_x[15731:15726] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15731:15726] * PIXEL_SIZE && v_count < i_worm_y[15731:15726] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2622 < i_size && h_count >= i_worm_x[15737:15732] * PIXEL_SIZE && h_count < i_worm_x[15737:15732] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15737:15732] * PIXEL_SIZE && v_count < i_worm_y[15737:15732] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2623 < i_size && h_count >= i_worm_x[15743:15738] * PIXEL_SIZE && h_count < i_worm_x[15743:15738] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15743:15738] * PIXEL_SIZE && v_count < i_worm_y[15743:15738] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2624 < i_size && h_count >= i_worm_x[15749:15744] * PIXEL_SIZE && h_count < i_worm_x[15749:15744] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15749:15744] * PIXEL_SIZE && v_count < i_worm_y[15749:15744] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2625 < i_size && h_count >= i_worm_x[15755:15750] * PIXEL_SIZE && h_count < i_worm_x[15755:15750] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15755:15750] * PIXEL_SIZE && v_count < i_worm_y[15755:15750] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2626 < i_size && h_count >= i_worm_x[15761:15756] * PIXEL_SIZE && h_count < i_worm_x[15761:15756] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15761:15756] * PIXEL_SIZE && v_count < i_worm_y[15761:15756] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2627 < i_size && h_count >= i_worm_x[15767:15762] * PIXEL_SIZE && h_count < i_worm_x[15767:15762] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15767:15762] * PIXEL_SIZE && v_count < i_worm_y[15767:15762] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2628 < i_size && h_count >= i_worm_x[15773:15768] * PIXEL_SIZE && h_count < i_worm_x[15773:15768] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15773:15768] * PIXEL_SIZE && v_count < i_worm_y[15773:15768] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2629 < i_size && h_count >= i_worm_x[15779:15774] * PIXEL_SIZE && h_count < i_worm_x[15779:15774] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15779:15774] * PIXEL_SIZE && v_count < i_worm_y[15779:15774] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2630 < i_size && h_count >= i_worm_x[15785:15780] * PIXEL_SIZE && h_count < i_worm_x[15785:15780] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15785:15780] * PIXEL_SIZE && v_count < i_worm_y[15785:15780] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2631 < i_size && h_count >= i_worm_x[15791:15786] * PIXEL_SIZE && h_count < i_worm_x[15791:15786] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15791:15786] * PIXEL_SIZE && v_count < i_worm_y[15791:15786] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2632 < i_size && h_count >= i_worm_x[15797:15792] * PIXEL_SIZE && h_count < i_worm_x[15797:15792] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15797:15792] * PIXEL_SIZE && v_count < i_worm_y[15797:15792] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2633 < i_size && h_count >= i_worm_x[15803:15798] * PIXEL_SIZE && h_count < i_worm_x[15803:15798] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15803:15798] * PIXEL_SIZE && v_count < i_worm_y[15803:15798] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2634 < i_size && h_count >= i_worm_x[15809:15804] * PIXEL_SIZE && h_count < i_worm_x[15809:15804] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15809:15804] * PIXEL_SIZE && v_count < i_worm_y[15809:15804] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2635 < i_size && h_count >= i_worm_x[15815:15810] * PIXEL_SIZE && h_count < i_worm_x[15815:15810] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15815:15810] * PIXEL_SIZE && v_count < i_worm_y[15815:15810] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2636 < i_size && h_count >= i_worm_x[15821:15816] * PIXEL_SIZE && h_count < i_worm_x[15821:15816] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15821:15816] * PIXEL_SIZE && v_count < i_worm_y[15821:15816] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2637 < i_size && h_count >= i_worm_x[15827:15822] * PIXEL_SIZE && h_count < i_worm_x[15827:15822] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15827:15822] * PIXEL_SIZE && v_count < i_worm_y[15827:15822] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2638 < i_size && h_count >= i_worm_x[15833:15828] * PIXEL_SIZE && h_count < i_worm_x[15833:15828] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15833:15828] * PIXEL_SIZE && v_count < i_worm_y[15833:15828] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2639 < i_size && h_count >= i_worm_x[15839:15834] * PIXEL_SIZE && h_count < i_worm_x[15839:15834] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15839:15834] * PIXEL_SIZE && v_count < i_worm_y[15839:15834] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2640 < i_size && h_count >= i_worm_x[15845:15840] * PIXEL_SIZE && h_count < i_worm_x[15845:15840] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15845:15840] * PIXEL_SIZE && v_count < i_worm_y[15845:15840] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2641 < i_size && h_count >= i_worm_x[15851:15846] * PIXEL_SIZE && h_count < i_worm_x[15851:15846] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15851:15846] * PIXEL_SIZE && v_count < i_worm_y[15851:15846] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2642 < i_size && h_count >= i_worm_x[15857:15852] * PIXEL_SIZE && h_count < i_worm_x[15857:15852] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15857:15852] * PIXEL_SIZE && v_count < i_worm_y[15857:15852] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2643 < i_size && h_count >= i_worm_x[15863:15858] * PIXEL_SIZE && h_count < i_worm_x[15863:15858] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15863:15858] * PIXEL_SIZE && v_count < i_worm_y[15863:15858] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2644 < i_size && h_count >= i_worm_x[15869:15864] * PIXEL_SIZE && h_count < i_worm_x[15869:15864] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15869:15864] * PIXEL_SIZE && v_count < i_worm_y[15869:15864] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2645 < i_size && h_count >= i_worm_x[15875:15870] * PIXEL_SIZE && h_count < i_worm_x[15875:15870] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15875:15870] * PIXEL_SIZE && v_count < i_worm_y[15875:15870] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2646 < i_size && h_count >= i_worm_x[15881:15876] * PIXEL_SIZE && h_count < i_worm_x[15881:15876] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15881:15876] * PIXEL_SIZE && v_count < i_worm_y[15881:15876] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2647 < i_size && h_count >= i_worm_x[15887:15882] * PIXEL_SIZE && h_count < i_worm_x[15887:15882] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15887:15882] * PIXEL_SIZE && v_count < i_worm_y[15887:15882] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2648 < i_size && h_count >= i_worm_x[15893:15888] * PIXEL_SIZE && h_count < i_worm_x[15893:15888] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15893:15888] * PIXEL_SIZE && v_count < i_worm_y[15893:15888] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2649 < i_size && h_count >= i_worm_x[15899:15894] * PIXEL_SIZE && h_count < i_worm_x[15899:15894] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15899:15894] * PIXEL_SIZE && v_count < i_worm_y[15899:15894] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2650 < i_size && h_count >= i_worm_x[15905:15900] * PIXEL_SIZE && h_count < i_worm_x[15905:15900] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15905:15900] * PIXEL_SIZE && v_count < i_worm_y[15905:15900] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2651 < i_size && h_count >= i_worm_x[15911:15906] * PIXEL_SIZE && h_count < i_worm_x[15911:15906] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15911:15906] * PIXEL_SIZE && v_count < i_worm_y[15911:15906] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2652 < i_size && h_count >= i_worm_x[15917:15912] * PIXEL_SIZE && h_count < i_worm_x[15917:15912] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15917:15912] * PIXEL_SIZE && v_count < i_worm_y[15917:15912] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2653 < i_size && h_count >= i_worm_x[15923:15918] * PIXEL_SIZE && h_count < i_worm_x[15923:15918] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15923:15918] * PIXEL_SIZE && v_count < i_worm_y[15923:15918] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2654 < i_size && h_count >= i_worm_x[15929:15924] * PIXEL_SIZE && h_count < i_worm_x[15929:15924] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15929:15924] * PIXEL_SIZE && v_count < i_worm_y[15929:15924] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2655 < i_size && h_count >= i_worm_x[15935:15930] * PIXEL_SIZE && h_count < i_worm_x[15935:15930] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15935:15930] * PIXEL_SIZE && v_count < i_worm_y[15935:15930] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2656 < i_size && h_count >= i_worm_x[15941:15936] * PIXEL_SIZE && h_count < i_worm_x[15941:15936] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15941:15936] * PIXEL_SIZE && v_count < i_worm_y[15941:15936] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2657 < i_size && h_count >= i_worm_x[15947:15942] * PIXEL_SIZE && h_count < i_worm_x[15947:15942] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15947:15942] * PIXEL_SIZE && v_count < i_worm_y[15947:15942] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2658 < i_size && h_count >= i_worm_x[15953:15948] * PIXEL_SIZE && h_count < i_worm_x[15953:15948] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15953:15948] * PIXEL_SIZE && v_count < i_worm_y[15953:15948] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2659 < i_size && h_count >= i_worm_x[15959:15954] * PIXEL_SIZE && h_count < i_worm_x[15959:15954] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15959:15954] * PIXEL_SIZE && v_count < i_worm_y[15959:15954] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2660 < i_size && h_count >= i_worm_x[15965:15960] * PIXEL_SIZE && h_count < i_worm_x[15965:15960] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15965:15960] * PIXEL_SIZE && v_count < i_worm_y[15965:15960] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2661 < i_size && h_count >= i_worm_x[15971:15966] * PIXEL_SIZE && h_count < i_worm_x[15971:15966] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15971:15966] * PIXEL_SIZE && v_count < i_worm_y[15971:15966] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2662 < i_size && h_count >= i_worm_x[15977:15972] * PIXEL_SIZE && h_count < i_worm_x[15977:15972] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15977:15972] * PIXEL_SIZE && v_count < i_worm_y[15977:15972] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2663 < i_size && h_count >= i_worm_x[15983:15978] * PIXEL_SIZE && h_count < i_worm_x[15983:15978] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15983:15978] * PIXEL_SIZE && v_count < i_worm_y[15983:15978] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2664 < i_size && h_count >= i_worm_x[15989:15984] * PIXEL_SIZE && h_count < i_worm_x[15989:15984] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15989:15984] * PIXEL_SIZE && v_count < i_worm_y[15989:15984] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2665 < i_size && h_count >= i_worm_x[15995:15990] * PIXEL_SIZE && h_count < i_worm_x[15995:15990] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[15995:15990] * PIXEL_SIZE && v_count < i_worm_y[15995:15990] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2666 < i_size && h_count >= i_worm_x[16001:15996] * PIXEL_SIZE && h_count < i_worm_x[16001:15996] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16001:15996] * PIXEL_SIZE && v_count < i_worm_y[16001:15996] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2667 < i_size && h_count >= i_worm_x[16007:16002] * PIXEL_SIZE && h_count < i_worm_x[16007:16002] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16007:16002] * PIXEL_SIZE && v_count < i_worm_y[16007:16002] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2668 < i_size && h_count >= i_worm_x[16013:16008] * PIXEL_SIZE && h_count < i_worm_x[16013:16008] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16013:16008] * PIXEL_SIZE && v_count < i_worm_y[16013:16008] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2669 < i_size && h_count >= i_worm_x[16019:16014] * PIXEL_SIZE && h_count < i_worm_x[16019:16014] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16019:16014] * PIXEL_SIZE && v_count < i_worm_y[16019:16014] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2670 < i_size && h_count >= i_worm_x[16025:16020] * PIXEL_SIZE && h_count < i_worm_x[16025:16020] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16025:16020] * PIXEL_SIZE && v_count < i_worm_y[16025:16020] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2671 < i_size && h_count >= i_worm_x[16031:16026] * PIXEL_SIZE && h_count < i_worm_x[16031:16026] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16031:16026] * PIXEL_SIZE && v_count < i_worm_y[16031:16026] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2672 < i_size && h_count >= i_worm_x[16037:16032] * PIXEL_SIZE && h_count < i_worm_x[16037:16032] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16037:16032] * PIXEL_SIZE && v_count < i_worm_y[16037:16032] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2673 < i_size && h_count >= i_worm_x[16043:16038] * PIXEL_SIZE && h_count < i_worm_x[16043:16038] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16043:16038] * PIXEL_SIZE && v_count < i_worm_y[16043:16038] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2674 < i_size && h_count >= i_worm_x[16049:16044] * PIXEL_SIZE && h_count < i_worm_x[16049:16044] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16049:16044] * PIXEL_SIZE && v_count < i_worm_y[16049:16044] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2675 < i_size && h_count >= i_worm_x[16055:16050] * PIXEL_SIZE && h_count < i_worm_x[16055:16050] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16055:16050] * PIXEL_SIZE && v_count < i_worm_y[16055:16050] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2676 < i_size && h_count >= i_worm_x[16061:16056] * PIXEL_SIZE && h_count < i_worm_x[16061:16056] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16061:16056] * PIXEL_SIZE && v_count < i_worm_y[16061:16056] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2677 < i_size && h_count >= i_worm_x[16067:16062] * PIXEL_SIZE && h_count < i_worm_x[16067:16062] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16067:16062] * PIXEL_SIZE && v_count < i_worm_y[16067:16062] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2678 < i_size && h_count >= i_worm_x[16073:16068] * PIXEL_SIZE && h_count < i_worm_x[16073:16068] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16073:16068] * PIXEL_SIZE && v_count < i_worm_y[16073:16068] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2679 < i_size && h_count >= i_worm_x[16079:16074] * PIXEL_SIZE && h_count < i_worm_x[16079:16074] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16079:16074] * PIXEL_SIZE && v_count < i_worm_y[16079:16074] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2680 < i_size && h_count >= i_worm_x[16085:16080] * PIXEL_SIZE && h_count < i_worm_x[16085:16080] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16085:16080] * PIXEL_SIZE && v_count < i_worm_y[16085:16080] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2681 < i_size && h_count >= i_worm_x[16091:16086] * PIXEL_SIZE && h_count < i_worm_x[16091:16086] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16091:16086] * PIXEL_SIZE && v_count < i_worm_y[16091:16086] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2682 < i_size && h_count >= i_worm_x[16097:16092] * PIXEL_SIZE && h_count < i_worm_x[16097:16092] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16097:16092] * PIXEL_SIZE && v_count < i_worm_y[16097:16092] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2683 < i_size && h_count >= i_worm_x[16103:16098] * PIXEL_SIZE && h_count < i_worm_x[16103:16098] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16103:16098] * PIXEL_SIZE && v_count < i_worm_y[16103:16098] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2684 < i_size && h_count >= i_worm_x[16109:16104] * PIXEL_SIZE && h_count < i_worm_x[16109:16104] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16109:16104] * PIXEL_SIZE && v_count < i_worm_y[16109:16104] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2685 < i_size && h_count >= i_worm_x[16115:16110] * PIXEL_SIZE && h_count < i_worm_x[16115:16110] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16115:16110] * PIXEL_SIZE && v_count < i_worm_y[16115:16110] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2686 < i_size && h_count >= i_worm_x[16121:16116] * PIXEL_SIZE && h_count < i_worm_x[16121:16116] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16121:16116] * PIXEL_SIZE && v_count < i_worm_y[16121:16116] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2687 < i_size && h_count >= i_worm_x[16127:16122] * PIXEL_SIZE && h_count < i_worm_x[16127:16122] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16127:16122] * PIXEL_SIZE && v_count < i_worm_y[16127:16122] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2688 < i_size && h_count >= i_worm_x[16133:16128] * PIXEL_SIZE && h_count < i_worm_x[16133:16128] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16133:16128] * PIXEL_SIZE && v_count < i_worm_y[16133:16128] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2689 < i_size && h_count >= i_worm_x[16139:16134] * PIXEL_SIZE && h_count < i_worm_x[16139:16134] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16139:16134] * PIXEL_SIZE && v_count < i_worm_y[16139:16134] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2690 < i_size && h_count >= i_worm_x[16145:16140] * PIXEL_SIZE && h_count < i_worm_x[16145:16140] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16145:16140] * PIXEL_SIZE && v_count < i_worm_y[16145:16140] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2691 < i_size && h_count >= i_worm_x[16151:16146] * PIXEL_SIZE && h_count < i_worm_x[16151:16146] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16151:16146] * PIXEL_SIZE && v_count < i_worm_y[16151:16146] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2692 < i_size && h_count >= i_worm_x[16157:16152] * PIXEL_SIZE && h_count < i_worm_x[16157:16152] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16157:16152] * PIXEL_SIZE && v_count < i_worm_y[16157:16152] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2693 < i_size && h_count >= i_worm_x[16163:16158] * PIXEL_SIZE && h_count < i_worm_x[16163:16158] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16163:16158] * PIXEL_SIZE && v_count < i_worm_y[16163:16158] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2694 < i_size && h_count >= i_worm_x[16169:16164] * PIXEL_SIZE && h_count < i_worm_x[16169:16164] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16169:16164] * PIXEL_SIZE && v_count < i_worm_y[16169:16164] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2695 < i_size && h_count >= i_worm_x[16175:16170] * PIXEL_SIZE && h_count < i_worm_x[16175:16170] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16175:16170] * PIXEL_SIZE && v_count < i_worm_y[16175:16170] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2696 < i_size && h_count >= i_worm_x[16181:16176] * PIXEL_SIZE && h_count < i_worm_x[16181:16176] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16181:16176] * PIXEL_SIZE && v_count < i_worm_y[16181:16176] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2697 < i_size && h_count >= i_worm_x[16187:16182] * PIXEL_SIZE && h_count < i_worm_x[16187:16182] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16187:16182] * PIXEL_SIZE && v_count < i_worm_y[16187:16182] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2698 < i_size && h_count >= i_worm_x[16193:16188] * PIXEL_SIZE && h_count < i_worm_x[16193:16188] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16193:16188] * PIXEL_SIZE && v_count < i_worm_y[16193:16188] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2699 < i_size && h_count >= i_worm_x[16199:16194] * PIXEL_SIZE && h_count < i_worm_x[16199:16194] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16199:16194] * PIXEL_SIZE && v_count < i_worm_y[16199:16194] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2700 < i_size && h_count >= i_worm_x[16205:16200] * PIXEL_SIZE && h_count < i_worm_x[16205:16200] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16205:16200] * PIXEL_SIZE && v_count < i_worm_y[16205:16200] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2701 < i_size && h_count >= i_worm_x[16211:16206] * PIXEL_SIZE && h_count < i_worm_x[16211:16206] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16211:16206] * PIXEL_SIZE && v_count < i_worm_y[16211:16206] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2702 < i_size && h_count >= i_worm_x[16217:16212] * PIXEL_SIZE && h_count < i_worm_x[16217:16212] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16217:16212] * PIXEL_SIZE && v_count < i_worm_y[16217:16212] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2703 < i_size && h_count >= i_worm_x[16223:16218] * PIXEL_SIZE && h_count < i_worm_x[16223:16218] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16223:16218] * PIXEL_SIZE && v_count < i_worm_y[16223:16218] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2704 < i_size && h_count >= i_worm_x[16229:16224] * PIXEL_SIZE && h_count < i_worm_x[16229:16224] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16229:16224] * PIXEL_SIZE && v_count < i_worm_y[16229:16224] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2705 < i_size && h_count >= i_worm_x[16235:16230] * PIXEL_SIZE && h_count < i_worm_x[16235:16230] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16235:16230] * PIXEL_SIZE && v_count < i_worm_y[16235:16230] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2706 < i_size && h_count >= i_worm_x[16241:16236] * PIXEL_SIZE && h_count < i_worm_x[16241:16236] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16241:16236] * PIXEL_SIZE && v_count < i_worm_y[16241:16236] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2707 < i_size && h_count >= i_worm_x[16247:16242] * PIXEL_SIZE && h_count < i_worm_x[16247:16242] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16247:16242] * PIXEL_SIZE && v_count < i_worm_y[16247:16242] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2708 < i_size && h_count >= i_worm_x[16253:16248] * PIXEL_SIZE && h_count < i_worm_x[16253:16248] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16253:16248] * PIXEL_SIZE && v_count < i_worm_y[16253:16248] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2709 < i_size && h_count >= i_worm_x[16259:16254] * PIXEL_SIZE && h_count < i_worm_x[16259:16254] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16259:16254] * PIXEL_SIZE && v_count < i_worm_y[16259:16254] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2710 < i_size && h_count >= i_worm_x[16265:16260] * PIXEL_SIZE && h_count < i_worm_x[16265:16260] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16265:16260] * PIXEL_SIZE && v_count < i_worm_y[16265:16260] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2711 < i_size && h_count >= i_worm_x[16271:16266] * PIXEL_SIZE && h_count < i_worm_x[16271:16266] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16271:16266] * PIXEL_SIZE && v_count < i_worm_y[16271:16266] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2712 < i_size && h_count >= i_worm_x[16277:16272] * PIXEL_SIZE && h_count < i_worm_x[16277:16272] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16277:16272] * PIXEL_SIZE && v_count < i_worm_y[16277:16272] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2713 < i_size && h_count >= i_worm_x[16283:16278] * PIXEL_SIZE && h_count < i_worm_x[16283:16278] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16283:16278] * PIXEL_SIZE && v_count < i_worm_y[16283:16278] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2714 < i_size && h_count >= i_worm_x[16289:16284] * PIXEL_SIZE && h_count < i_worm_x[16289:16284] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16289:16284] * PIXEL_SIZE && v_count < i_worm_y[16289:16284] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2715 < i_size && h_count >= i_worm_x[16295:16290] * PIXEL_SIZE && h_count < i_worm_x[16295:16290] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16295:16290] * PIXEL_SIZE && v_count < i_worm_y[16295:16290] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2716 < i_size && h_count >= i_worm_x[16301:16296] * PIXEL_SIZE && h_count < i_worm_x[16301:16296] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16301:16296] * PIXEL_SIZE && v_count < i_worm_y[16301:16296] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2717 < i_size && h_count >= i_worm_x[16307:16302] * PIXEL_SIZE && h_count < i_worm_x[16307:16302] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16307:16302] * PIXEL_SIZE && v_count < i_worm_y[16307:16302] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2718 < i_size && h_count >= i_worm_x[16313:16308] * PIXEL_SIZE && h_count < i_worm_x[16313:16308] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16313:16308] * PIXEL_SIZE && v_count < i_worm_y[16313:16308] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2719 < i_size && h_count >= i_worm_x[16319:16314] * PIXEL_SIZE && h_count < i_worm_x[16319:16314] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16319:16314] * PIXEL_SIZE && v_count < i_worm_y[16319:16314] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2720 < i_size && h_count >= i_worm_x[16325:16320] * PIXEL_SIZE && h_count < i_worm_x[16325:16320] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16325:16320] * PIXEL_SIZE && v_count < i_worm_y[16325:16320] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2721 < i_size && h_count >= i_worm_x[16331:16326] * PIXEL_SIZE && h_count < i_worm_x[16331:16326] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16331:16326] * PIXEL_SIZE && v_count < i_worm_y[16331:16326] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2722 < i_size && h_count >= i_worm_x[16337:16332] * PIXEL_SIZE && h_count < i_worm_x[16337:16332] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16337:16332] * PIXEL_SIZE && v_count < i_worm_y[16337:16332] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2723 < i_size && h_count >= i_worm_x[16343:16338] * PIXEL_SIZE && h_count < i_worm_x[16343:16338] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16343:16338] * PIXEL_SIZE && v_count < i_worm_y[16343:16338] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2724 < i_size && h_count >= i_worm_x[16349:16344] * PIXEL_SIZE && h_count < i_worm_x[16349:16344] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16349:16344] * PIXEL_SIZE && v_count < i_worm_y[16349:16344] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2725 < i_size && h_count >= i_worm_x[16355:16350] * PIXEL_SIZE && h_count < i_worm_x[16355:16350] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16355:16350] * PIXEL_SIZE && v_count < i_worm_y[16355:16350] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2726 < i_size && h_count >= i_worm_x[16361:16356] * PIXEL_SIZE && h_count < i_worm_x[16361:16356] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16361:16356] * PIXEL_SIZE && v_count < i_worm_y[16361:16356] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2727 < i_size && h_count >= i_worm_x[16367:16362] * PIXEL_SIZE && h_count < i_worm_x[16367:16362] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16367:16362] * PIXEL_SIZE && v_count < i_worm_y[16367:16362] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2728 < i_size && h_count >= i_worm_x[16373:16368] * PIXEL_SIZE && h_count < i_worm_x[16373:16368] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16373:16368] * PIXEL_SIZE && v_count < i_worm_y[16373:16368] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2729 < i_size && h_count >= i_worm_x[16379:16374] * PIXEL_SIZE && h_count < i_worm_x[16379:16374] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16379:16374] * PIXEL_SIZE && v_count < i_worm_y[16379:16374] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2730 < i_size && h_count >= i_worm_x[16385:16380] * PIXEL_SIZE && h_count < i_worm_x[16385:16380] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16385:16380] * PIXEL_SIZE && v_count < i_worm_y[16385:16380] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2731 < i_size && h_count >= i_worm_x[16391:16386] * PIXEL_SIZE && h_count < i_worm_x[16391:16386] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16391:16386] * PIXEL_SIZE && v_count < i_worm_y[16391:16386] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2732 < i_size && h_count >= i_worm_x[16397:16392] * PIXEL_SIZE && h_count < i_worm_x[16397:16392] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16397:16392] * PIXEL_SIZE && v_count < i_worm_y[16397:16392] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2733 < i_size && h_count >= i_worm_x[16403:16398] * PIXEL_SIZE && h_count < i_worm_x[16403:16398] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16403:16398] * PIXEL_SIZE && v_count < i_worm_y[16403:16398] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2734 < i_size && h_count >= i_worm_x[16409:16404] * PIXEL_SIZE && h_count < i_worm_x[16409:16404] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16409:16404] * PIXEL_SIZE && v_count < i_worm_y[16409:16404] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2735 < i_size && h_count >= i_worm_x[16415:16410] * PIXEL_SIZE && h_count < i_worm_x[16415:16410] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16415:16410] * PIXEL_SIZE && v_count < i_worm_y[16415:16410] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2736 < i_size && h_count >= i_worm_x[16421:16416] * PIXEL_SIZE && h_count < i_worm_x[16421:16416] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16421:16416] * PIXEL_SIZE && v_count < i_worm_y[16421:16416] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2737 < i_size && h_count >= i_worm_x[16427:16422] * PIXEL_SIZE && h_count < i_worm_x[16427:16422] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16427:16422] * PIXEL_SIZE && v_count < i_worm_y[16427:16422] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2738 < i_size && h_count >= i_worm_x[16433:16428] * PIXEL_SIZE && h_count < i_worm_x[16433:16428] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16433:16428] * PIXEL_SIZE && v_count < i_worm_y[16433:16428] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2739 < i_size && h_count >= i_worm_x[16439:16434] * PIXEL_SIZE && h_count < i_worm_x[16439:16434] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16439:16434] * PIXEL_SIZE && v_count < i_worm_y[16439:16434] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2740 < i_size && h_count >= i_worm_x[16445:16440] * PIXEL_SIZE && h_count < i_worm_x[16445:16440] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16445:16440] * PIXEL_SIZE && v_count < i_worm_y[16445:16440] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2741 < i_size && h_count >= i_worm_x[16451:16446] * PIXEL_SIZE && h_count < i_worm_x[16451:16446] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16451:16446] * PIXEL_SIZE && v_count < i_worm_y[16451:16446] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2742 < i_size && h_count >= i_worm_x[16457:16452] * PIXEL_SIZE && h_count < i_worm_x[16457:16452] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16457:16452] * PIXEL_SIZE && v_count < i_worm_y[16457:16452] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2743 < i_size && h_count >= i_worm_x[16463:16458] * PIXEL_SIZE && h_count < i_worm_x[16463:16458] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16463:16458] * PIXEL_SIZE && v_count < i_worm_y[16463:16458] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2744 < i_size && h_count >= i_worm_x[16469:16464] * PIXEL_SIZE && h_count < i_worm_x[16469:16464] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16469:16464] * PIXEL_SIZE && v_count < i_worm_y[16469:16464] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2745 < i_size && h_count >= i_worm_x[16475:16470] * PIXEL_SIZE && h_count < i_worm_x[16475:16470] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16475:16470] * PIXEL_SIZE && v_count < i_worm_y[16475:16470] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2746 < i_size && h_count >= i_worm_x[16481:16476] * PIXEL_SIZE && h_count < i_worm_x[16481:16476] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16481:16476] * PIXEL_SIZE && v_count < i_worm_y[16481:16476] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2747 < i_size && h_count >= i_worm_x[16487:16482] * PIXEL_SIZE && h_count < i_worm_x[16487:16482] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16487:16482] * PIXEL_SIZE && v_count < i_worm_y[16487:16482] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2748 < i_size && h_count >= i_worm_x[16493:16488] * PIXEL_SIZE && h_count < i_worm_x[16493:16488] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16493:16488] * PIXEL_SIZE && v_count < i_worm_y[16493:16488] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2749 < i_size && h_count >= i_worm_x[16499:16494] * PIXEL_SIZE && h_count < i_worm_x[16499:16494] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16499:16494] * PIXEL_SIZE && v_count < i_worm_y[16499:16494] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2750 < i_size && h_count >= i_worm_x[16505:16500] * PIXEL_SIZE && h_count < i_worm_x[16505:16500] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16505:16500] * PIXEL_SIZE && v_count < i_worm_y[16505:16500] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2751 < i_size && h_count >= i_worm_x[16511:16506] * PIXEL_SIZE && h_count < i_worm_x[16511:16506] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16511:16506] * PIXEL_SIZE && v_count < i_worm_y[16511:16506] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2752 < i_size && h_count >= i_worm_x[16517:16512] * PIXEL_SIZE && h_count < i_worm_x[16517:16512] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16517:16512] * PIXEL_SIZE && v_count < i_worm_y[16517:16512] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2753 < i_size && h_count >= i_worm_x[16523:16518] * PIXEL_SIZE && h_count < i_worm_x[16523:16518] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16523:16518] * PIXEL_SIZE && v_count < i_worm_y[16523:16518] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2754 < i_size && h_count >= i_worm_x[16529:16524] * PIXEL_SIZE && h_count < i_worm_x[16529:16524] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16529:16524] * PIXEL_SIZE && v_count < i_worm_y[16529:16524] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2755 < i_size && h_count >= i_worm_x[16535:16530] * PIXEL_SIZE && h_count < i_worm_x[16535:16530] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16535:16530] * PIXEL_SIZE && v_count < i_worm_y[16535:16530] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2756 < i_size && h_count >= i_worm_x[16541:16536] * PIXEL_SIZE && h_count < i_worm_x[16541:16536] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16541:16536] * PIXEL_SIZE && v_count < i_worm_y[16541:16536] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2757 < i_size && h_count >= i_worm_x[16547:16542] * PIXEL_SIZE && h_count < i_worm_x[16547:16542] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16547:16542] * PIXEL_SIZE && v_count < i_worm_y[16547:16542] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2758 < i_size && h_count >= i_worm_x[16553:16548] * PIXEL_SIZE && h_count < i_worm_x[16553:16548] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16553:16548] * PIXEL_SIZE && v_count < i_worm_y[16553:16548] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2759 < i_size && h_count >= i_worm_x[16559:16554] * PIXEL_SIZE && h_count < i_worm_x[16559:16554] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16559:16554] * PIXEL_SIZE && v_count < i_worm_y[16559:16554] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2760 < i_size && h_count >= i_worm_x[16565:16560] * PIXEL_SIZE && h_count < i_worm_x[16565:16560] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16565:16560] * PIXEL_SIZE && v_count < i_worm_y[16565:16560] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2761 < i_size && h_count >= i_worm_x[16571:16566] * PIXEL_SIZE && h_count < i_worm_x[16571:16566] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16571:16566] * PIXEL_SIZE && v_count < i_worm_y[16571:16566] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2762 < i_size && h_count >= i_worm_x[16577:16572] * PIXEL_SIZE && h_count < i_worm_x[16577:16572] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16577:16572] * PIXEL_SIZE && v_count < i_worm_y[16577:16572] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2763 < i_size && h_count >= i_worm_x[16583:16578] * PIXEL_SIZE && h_count < i_worm_x[16583:16578] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16583:16578] * PIXEL_SIZE && v_count < i_worm_y[16583:16578] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2764 < i_size && h_count >= i_worm_x[16589:16584] * PIXEL_SIZE && h_count < i_worm_x[16589:16584] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16589:16584] * PIXEL_SIZE && v_count < i_worm_y[16589:16584] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2765 < i_size && h_count >= i_worm_x[16595:16590] * PIXEL_SIZE && h_count < i_worm_x[16595:16590] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16595:16590] * PIXEL_SIZE && v_count < i_worm_y[16595:16590] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2766 < i_size && h_count >= i_worm_x[16601:16596] * PIXEL_SIZE && h_count < i_worm_x[16601:16596] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16601:16596] * PIXEL_SIZE && v_count < i_worm_y[16601:16596] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2767 < i_size && h_count >= i_worm_x[16607:16602] * PIXEL_SIZE && h_count < i_worm_x[16607:16602] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16607:16602] * PIXEL_SIZE && v_count < i_worm_y[16607:16602] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2768 < i_size && h_count >= i_worm_x[16613:16608] * PIXEL_SIZE && h_count < i_worm_x[16613:16608] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16613:16608] * PIXEL_SIZE && v_count < i_worm_y[16613:16608] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2769 < i_size && h_count >= i_worm_x[16619:16614] * PIXEL_SIZE && h_count < i_worm_x[16619:16614] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16619:16614] * PIXEL_SIZE && v_count < i_worm_y[16619:16614] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2770 < i_size && h_count >= i_worm_x[16625:16620] * PIXEL_SIZE && h_count < i_worm_x[16625:16620] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16625:16620] * PIXEL_SIZE && v_count < i_worm_y[16625:16620] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2771 < i_size && h_count >= i_worm_x[16631:16626] * PIXEL_SIZE && h_count < i_worm_x[16631:16626] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16631:16626] * PIXEL_SIZE && v_count < i_worm_y[16631:16626] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2772 < i_size && h_count >= i_worm_x[16637:16632] * PIXEL_SIZE && h_count < i_worm_x[16637:16632] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16637:16632] * PIXEL_SIZE && v_count < i_worm_y[16637:16632] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2773 < i_size && h_count >= i_worm_x[16643:16638] * PIXEL_SIZE && h_count < i_worm_x[16643:16638] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16643:16638] * PIXEL_SIZE && v_count < i_worm_y[16643:16638] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2774 < i_size && h_count >= i_worm_x[16649:16644] * PIXEL_SIZE && h_count < i_worm_x[16649:16644] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16649:16644] * PIXEL_SIZE && v_count < i_worm_y[16649:16644] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2775 < i_size && h_count >= i_worm_x[16655:16650] * PIXEL_SIZE && h_count < i_worm_x[16655:16650] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16655:16650] * PIXEL_SIZE && v_count < i_worm_y[16655:16650] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2776 < i_size && h_count >= i_worm_x[16661:16656] * PIXEL_SIZE && h_count < i_worm_x[16661:16656] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16661:16656] * PIXEL_SIZE && v_count < i_worm_y[16661:16656] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2777 < i_size && h_count >= i_worm_x[16667:16662] * PIXEL_SIZE && h_count < i_worm_x[16667:16662] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16667:16662] * PIXEL_SIZE && v_count < i_worm_y[16667:16662] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2778 < i_size && h_count >= i_worm_x[16673:16668] * PIXEL_SIZE && h_count < i_worm_x[16673:16668] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16673:16668] * PIXEL_SIZE && v_count < i_worm_y[16673:16668] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2779 < i_size && h_count >= i_worm_x[16679:16674] * PIXEL_SIZE && h_count < i_worm_x[16679:16674] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16679:16674] * PIXEL_SIZE && v_count < i_worm_y[16679:16674] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2780 < i_size && h_count >= i_worm_x[16685:16680] * PIXEL_SIZE && h_count < i_worm_x[16685:16680] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16685:16680] * PIXEL_SIZE && v_count < i_worm_y[16685:16680] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2781 < i_size && h_count >= i_worm_x[16691:16686] * PIXEL_SIZE && h_count < i_worm_x[16691:16686] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16691:16686] * PIXEL_SIZE && v_count < i_worm_y[16691:16686] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2782 < i_size && h_count >= i_worm_x[16697:16692] * PIXEL_SIZE && h_count < i_worm_x[16697:16692] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16697:16692] * PIXEL_SIZE && v_count < i_worm_y[16697:16692] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2783 < i_size && h_count >= i_worm_x[16703:16698] * PIXEL_SIZE && h_count < i_worm_x[16703:16698] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16703:16698] * PIXEL_SIZE && v_count < i_worm_y[16703:16698] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2784 < i_size && h_count >= i_worm_x[16709:16704] * PIXEL_SIZE && h_count < i_worm_x[16709:16704] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16709:16704] * PIXEL_SIZE && v_count < i_worm_y[16709:16704] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2785 < i_size && h_count >= i_worm_x[16715:16710] * PIXEL_SIZE && h_count < i_worm_x[16715:16710] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16715:16710] * PIXEL_SIZE && v_count < i_worm_y[16715:16710] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2786 < i_size && h_count >= i_worm_x[16721:16716] * PIXEL_SIZE && h_count < i_worm_x[16721:16716] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16721:16716] * PIXEL_SIZE && v_count < i_worm_y[16721:16716] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2787 < i_size && h_count >= i_worm_x[16727:16722] * PIXEL_SIZE && h_count < i_worm_x[16727:16722] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16727:16722] * PIXEL_SIZE && v_count < i_worm_y[16727:16722] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2788 < i_size && h_count >= i_worm_x[16733:16728] * PIXEL_SIZE && h_count < i_worm_x[16733:16728] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16733:16728] * PIXEL_SIZE && v_count < i_worm_y[16733:16728] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2789 < i_size && h_count >= i_worm_x[16739:16734] * PIXEL_SIZE && h_count < i_worm_x[16739:16734] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16739:16734] * PIXEL_SIZE && v_count < i_worm_y[16739:16734] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2790 < i_size && h_count >= i_worm_x[16745:16740] * PIXEL_SIZE && h_count < i_worm_x[16745:16740] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16745:16740] * PIXEL_SIZE && v_count < i_worm_y[16745:16740] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2791 < i_size && h_count >= i_worm_x[16751:16746] * PIXEL_SIZE && h_count < i_worm_x[16751:16746] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16751:16746] * PIXEL_SIZE && v_count < i_worm_y[16751:16746] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2792 < i_size && h_count >= i_worm_x[16757:16752] * PIXEL_SIZE && h_count < i_worm_x[16757:16752] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16757:16752] * PIXEL_SIZE && v_count < i_worm_y[16757:16752] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2793 < i_size && h_count >= i_worm_x[16763:16758] * PIXEL_SIZE && h_count < i_worm_x[16763:16758] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16763:16758] * PIXEL_SIZE && v_count < i_worm_y[16763:16758] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2794 < i_size && h_count >= i_worm_x[16769:16764] * PIXEL_SIZE && h_count < i_worm_x[16769:16764] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16769:16764] * PIXEL_SIZE && v_count < i_worm_y[16769:16764] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2795 < i_size && h_count >= i_worm_x[16775:16770] * PIXEL_SIZE && h_count < i_worm_x[16775:16770] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16775:16770] * PIXEL_SIZE && v_count < i_worm_y[16775:16770] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2796 < i_size && h_count >= i_worm_x[16781:16776] * PIXEL_SIZE && h_count < i_worm_x[16781:16776] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16781:16776] * PIXEL_SIZE && v_count < i_worm_y[16781:16776] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2797 < i_size && h_count >= i_worm_x[16787:16782] * PIXEL_SIZE && h_count < i_worm_x[16787:16782] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16787:16782] * PIXEL_SIZE && v_count < i_worm_y[16787:16782] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2798 < i_size && h_count >= i_worm_x[16793:16788] * PIXEL_SIZE && h_count < i_worm_x[16793:16788] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16793:16788] * PIXEL_SIZE && v_count < i_worm_y[16793:16788] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2799 < i_size && h_count >= i_worm_x[16799:16794] * PIXEL_SIZE && h_count < i_worm_x[16799:16794] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16799:16794] * PIXEL_SIZE && v_count < i_worm_y[16799:16794] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2800 < i_size && h_count >= i_worm_x[16805:16800] * PIXEL_SIZE && h_count < i_worm_x[16805:16800] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16805:16800] * PIXEL_SIZE && v_count < i_worm_y[16805:16800] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2801 < i_size && h_count >= i_worm_x[16811:16806] * PIXEL_SIZE && h_count < i_worm_x[16811:16806] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16811:16806] * PIXEL_SIZE && v_count < i_worm_y[16811:16806] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2802 < i_size && h_count >= i_worm_x[16817:16812] * PIXEL_SIZE && h_count < i_worm_x[16817:16812] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16817:16812] * PIXEL_SIZE && v_count < i_worm_y[16817:16812] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2803 < i_size && h_count >= i_worm_x[16823:16818] * PIXEL_SIZE && h_count < i_worm_x[16823:16818] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16823:16818] * PIXEL_SIZE && v_count < i_worm_y[16823:16818] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2804 < i_size && h_count >= i_worm_x[16829:16824] * PIXEL_SIZE && h_count < i_worm_x[16829:16824] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16829:16824] * PIXEL_SIZE && v_count < i_worm_y[16829:16824] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2805 < i_size && h_count >= i_worm_x[16835:16830] * PIXEL_SIZE && h_count < i_worm_x[16835:16830] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16835:16830] * PIXEL_SIZE && v_count < i_worm_y[16835:16830] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2806 < i_size && h_count >= i_worm_x[16841:16836] * PIXEL_SIZE && h_count < i_worm_x[16841:16836] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16841:16836] * PIXEL_SIZE && v_count < i_worm_y[16841:16836] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2807 < i_size && h_count >= i_worm_x[16847:16842] * PIXEL_SIZE && h_count < i_worm_x[16847:16842] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16847:16842] * PIXEL_SIZE && v_count < i_worm_y[16847:16842] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2808 < i_size && h_count >= i_worm_x[16853:16848] * PIXEL_SIZE && h_count < i_worm_x[16853:16848] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16853:16848] * PIXEL_SIZE && v_count < i_worm_y[16853:16848] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2809 < i_size && h_count >= i_worm_x[16859:16854] * PIXEL_SIZE && h_count < i_worm_x[16859:16854] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16859:16854] * PIXEL_SIZE && v_count < i_worm_y[16859:16854] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2810 < i_size && h_count >= i_worm_x[16865:16860] * PIXEL_SIZE && h_count < i_worm_x[16865:16860] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16865:16860] * PIXEL_SIZE && v_count < i_worm_y[16865:16860] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2811 < i_size && h_count >= i_worm_x[16871:16866] * PIXEL_SIZE && h_count < i_worm_x[16871:16866] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16871:16866] * PIXEL_SIZE && v_count < i_worm_y[16871:16866] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2812 < i_size && h_count >= i_worm_x[16877:16872] * PIXEL_SIZE && h_count < i_worm_x[16877:16872] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16877:16872] * PIXEL_SIZE && v_count < i_worm_y[16877:16872] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2813 < i_size && h_count >= i_worm_x[16883:16878] * PIXEL_SIZE && h_count < i_worm_x[16883:16878] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16883:16878] * PIXEL_SIZE && v_count < i_worm_y[16883:16878] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2814 < i_size && h_count >= i_worm_x[16889:16884] * PIXEL_SIZE && h_count < i_worm_x[16889:16884] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16889:16884] * PIXEL_SIZE && v_count < i_worm_y[16889:16884] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2815 < i_size && h_count >= i_worm_x[16895:16890] * PIXEL_SIZE && h_count < i_worm_x[16895:16890] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16895:16890] * PIXEL_SIZE && v_count < i_worm_y[16895:16890] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2816 < i_size && h_count >= i_worm_x[16901:16896] * PIXEL_SIZE && h_count < i_worm_x[16901:16896] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16901:16896] * PIXEL_SIZE && v_count < i_worm_y[16901:16896] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2817 < i_size && h_count >= i_worm_x[16907:16902] * PIXEL_SIZE && h_count < i_worm_x[16907:16902] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16907:16902] * PIXEL_SIZE && v_count < i_worm_y[16907:16902] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2818 < i_size && h_count >= i_worm_x[16913:16908] * PIXEL_SIZE && h_count < i_worm_x[16913:16908] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16913:16908] * PIXEL_SIZE && v_count < i_worm_y[16913:16908] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2819 < i_size && h_count >= i_worm_x[16919:16914] * PIXEL_SIZE && h_count < i_worm_x[16919:16914] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16919:16914] * PIXEL_SIZE && v_count < i_worm_y[16919:16914] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2820 < i_size && h_count >= i_worm_x[16925:16920] * PIXEL_SIZE && h_count < i_worm_x[16925:16920] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16925:16920] * PIXEL_SIZE && v_count < i_worm_y[16925:16920] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2821 < i_size && h_count >= i_worm_x[16931:16926] * PIXEL_SIZE && h_count < i_worm_x[16931:16926] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16931:16926] * PIXEL_SIZE && v_count < i_worm_y[16931:16926] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2822 < i_size && h_count >= i_worm_x[16937:16932] * PIXEL_SIZE && h_count < i_worm_x[16937:16932] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16937:16932] * PIXEL_SIZE && v_count < i_worm_y[16937:16932] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2823 < i_size && h_count >= i_worm_x[16943:16938] * PIXEL_SIZE && h_count < i_worm_x[16943:16938] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16943:16938] * PIXEL_SIZE && v_count < i_worm_y[16943:16938] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2824 < i_size && h_count >= i_worm_x[16949:16944] * PIXEL_SIZE && h_count < i_worm_x[16949:16944] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16949:16944] * PIXEL_SIZE && v_count < i_worm_y[16949:16944] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2825 < i_size && h_count >= i_worm_x[16955:16950] * PIXEL_SIZE && h_count < i_worm_x[16955:16950] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16955:16950] * PIXEL_SIZE && v_count < i_worm_y[16955:16950] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2826 < i_size && h_count >= i_worm_x[16961:16956] * PIXEL_SIZE && h_count < i_worm_x[16961:16956] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16961:16956] * PIXEL_SIZE && v_count < i_worm_y[16961:16956] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2827 < i_size && h_count >= i_worm_x[16967:16962] * PIXEL_SIZE && h_count < i_worm_x[16967:16962] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16967:16962] * PIXEL_SIZE && v_count < i_worm_y[16967:16962] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2828 < i_size && h_count >= i_worm_x[16973:16968] * PIXEL_SIZE && h_count < i_worm_x[16973:16968] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16973:16968] * PIXEL_SIZE && v_count < i_worm_y[16973:16968] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2829 < i_size && h_count >= i_worm_x[16979:16974] * PIXEL_SIZE && h_count < i_worm_x[16979:16974] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16979:16974] * PIXEL_SIZE && v_count < i_worm_y[16979:16974] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2830 < i_size && h_count >= i_worm_x[16985:16980] * PIXEL_SIZE && h_count < i_worm_x[16985:16980] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16985:16980] * PIXEL_SIZE && v_count < i_worm_y[16985:16980] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2831 < i_size && h_count >= i_worm_x[16991:16986] * PIXEL_SIZE && h_count < i_worm_x[16991:16986] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16991:16986] * PIXEL_SIZE && v_count < i_worm_y[16991:16986] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2832 < i_size && h_count >= i_worm_x[16997:16992] * PIXEL_SIZE && h_count < i_worm_x[16997:16992] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[16997:16992] * PIXEL_SIZE && v_count < i_worm_y[16997:16992] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2833 < i_size && h_count >= i_worm_x[17003:16998] * PIXEL_SIZE && h_count < i_worm_x[17003:16998] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17003:16998] * PIXEL_SIZE && v_count < i_worm_y[17003:16998] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2834 < i_size && h_count >= i_worm_x[17009:17004] * PIXEL_SIZE && h_count < i_worm_x[17009:17004] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17009:17004] * PIXEL_SIZE && v_count < i_worm_y[17009:17004] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2835 < i_size && h_count >= i_worm_x[17015:17010] * PIXEL_SIZE && h_count < i_worm_x[17015:17010] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17015:17010] * PIXEL_SIZE && v_count < i_worm_y[17015:17010] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2836 < i_size && h_count >= i_worm_x[17021:17016] * PIXEL_SIZE && h_count < i_worm_x[17021:17016] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17021:17016] * PIXEL_SIZE && v_count < i_worm_y[17021:17016] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2837 < i_size && h_count >= i_worm_x[17027:17022] * PIXEL_SIZE && h_count < i_worm_x[17027:17022] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17027:17022] * PIXEL_SIZE && v_count < i_worm_y[17027:17022] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2838 < i_size && h_count >= i_worm_x[17033:17028] * PIXEL_SIZE && h_count < i_worm_x[17033:17028] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17033:17028] * PIXEL_SIZE && v_count < i_worm_y[17033:17028] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2839 < i_size && h_count >= i_worm_x[17039:17034] * PIXEL_SIZE && h_count < i_worm_x[17039:17034] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17039:17034] * PIXEL_SIZE && v_count < i_worm_y[17039:17034] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2840 < i_size && h_count >= i_worm_x[17045:17040] * PIXEL_SIZE && h_count < i_worm_x[17045:17040] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17045:17040] * PIXEL_SIZE && v_count < i_worm_y[17045:17040] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2841 < i_size && h_count >= i_worm_x[17051:17046] * PIXEL_SIZE && h_count < i_worm_x[17051:17046] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17051:17046] * PIXEL_SIZE && v_count < i_worm_y[17051:17046] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2842 < i_size && h_count >= i_worm_x[17057:17052] * PIXEL_SIZE && h_count < i_worm_x[17057:17052] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17057:17052] * PIXEL_SIZE && v_count < i_worm_y[17057:17052] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2843 < i_size && h_count >= i_worm_x[17063:17058] * PIXEL_SIZE && h_count < i_worm_x[17063:17058] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17063:17058] * PIXEL_SIZE && v_count < i_worm_y[17063:17058] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2844 < i_size && h_count >= i_worm_x[17069:17064] * PIXEL_SIZE && h_count < i_worm_x[17069:17064] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17069:17064] * PIXEL_SIZE && v_count < i_worm_y[17069:17064] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2845 < i_size && h_count >= i_worm_x[17075:17070] * PIXEL_SIZE && h_count < i_worm_x[17075:17070] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17075:17070] * PIXEL_SIZE && v_count < i_worm_y[17075:17070] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2846 < i_size && h_count >= i_worm_x[17081:17076] * PIXEL_SIZE && h_count < i_worm_x[17081:17076] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17081:17076] * PIXEL_SIZE && v_count < i_worm_y[17081:17076] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2847 < i_size && h_count >= i_worm_x[17087:17082] * PIXEL_SIZE && h_count < i_worm_x[17087:17082] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17087:17082] * PIXEL_SIZE && v_count < i_worm_y[17087:17082] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2848 < i_size && h_count >= i_worm_x[17093:17088] * PIXEL_SIZE && h_count < i_worm_x[17093:17088] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17093:17088] * PIXEL_SIZE && v_count < i_worm_y[17093:17088] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2849 < i_size && h_count >= i_worm_x[17099:17094] * PIXEL_SIZE && h_count < i_worm_x[17099:17094] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17099:17094] * PIXEL_SIZE && v_count < i_worm_y[17099:17094] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2850 < i_size && h_count >= i_worm_x[17105:17100] * PIXEL_SIZE && h_count < i_worm_x[17105:17100] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17105:17100] * PIXEL_SIZE && v_count < i_worm_y[17105:17100] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2851 < i_size && h_count >= i_worm_x[17111:17106] * PIXEL_SIZE && h_count < i_worm_x[17111:17106] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17111:17106] * PIXEL_SIZE && v_count < i_worm_y[17111:17106] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2852 < i_size && h_count >= i_worm_x[17117:17112] * PIXEL_SIZE && h_count < i_worm_x[17117:17112] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17117:17112] * PIXEL_SIZE && v_count < i_worm_y[17117:17112] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2853 < i_size && h_count >= i_worm_x[17123:17118] * PIXEL_SIZE && h_count < i_worm_x[17123:17118] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17123:17118] * PIXEL_SIZE && v_count < i_worm_y[17123:17118] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2854 < i_size && h_count >= i_worm_x[17129:17124] * PIXEL_SIZE && h_count < i_worm_x[17129:17124] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17129:17124] * PIXEL_SIZE && v_count < i_worm_y[17129:17124] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2855 < i_size && h_count >= i_worm_x[17135:17130] * PIXEL_SIZE && h_count < i_worm_x[17135:17130] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17135:17130] * PIXEL_SIZE && v_count < i_worm_y[17135:17130] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2856 < i_size && h_count >= i_worm_x[17141:17136] * PIXEL_SIZE && h_count < i_worm_x[17141:17136] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17141:17136] * PIXEL_SIZE && v_count < i_worm_y[17141:17136] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2857 < i_size && h_count >= i_worm_x[17147:17142] * PIXEL_SIZE && h_count < i_worm_x[17147:17142] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17147:17142] * PIXEL_SIZE && v_count < i_worm_y[17147:17142] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2858 < i_size && h_count >= i_worm_x[17153:17148] * PIXEL_SIZE && h_count < i_worm_x[17153:17148] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17153:17148] * PIXEL_SIZE && v_count < i_worm_y[17153:17148] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2859 < i_size && h_count >= i_worm_x[17159:17154] * PIXEL_SIZE && h_count < i_worm_x[17159:17154] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17159:17154] * PIXEL_SIZE && v_count < i_worm_y[17159:17154] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2860 < i_size && h_count >= i_worm_x[17165:17160] * PIXEL_SIZE && h_count < i_worm_x[17165:17160] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17165:17160] * PIXEL_SIZE && v_count < i_worm_y[17165:17160] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2861 < i_size && h_count >= i_worm_x[17171:17166] * PIXEL_SIZE && h_count < i_worm_x[17171:17166] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17171:17166] * PIXEL_SIZE && v_count < i_worm_y[17171:17166] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2862 < i_size && h_count >= i_worm_x[17177:17172] * PIXEL_SIZE && h_count < i_worm_x[17177:17172] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17177:17172] * PIXEL_SIZE && v_count < i_worm_y[17177:17172] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2863 < i_size && h_count >= i_worm_x[17183:17178] * PIXEL_SIZE && h_count < i_worm_x[17183:17178] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17183:17178] * PIXEL_SIZE && v_count < i_worm_y[17183:17178] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2864 < i_size && h_count >= i_worm_x[17189:17184] * PIXEL_SIZE && h_count < i_worm_x[17189:17184] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17189:17184] * PIXEL_SIZE && v_count < i_worm_y[17189:17184] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2865 < i_size && h_count >= i_worm_x[17195:17190] * PIXEL_SIZE && h_count < i_worm_x[17195:17190] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17195:17190] * PIXEL_SIZE && v_count < i_worm_y[17195:17190] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2866 < i_size && h_count >= i_worm_x[17201:17196] * PIXEL_SIZE && h_count < i_worm_x[17201:17196] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17201:17196] * PIXEL_SIZE && v_count < i_worm_y[17201:17196] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2867 < i_size && h_count >= i_worm_x[17207:17202] * PIXEL_SIZE && h_count < i_worm_x[17207:17202] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17207:17202] * PIXEL_SIZE && v_count < i_worm_y[17207:17202] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2868 < i_size && h_count >= i_worm_x[17213:17208] * PIXEL_SIZE && h_count < i_worm_x[17213:17208] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17213:17208] * PIXEL_SIZE && v_count < i_worm_y[17213:17208] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2869 < i_size && h_count >= i_worm_x[17219:17214] * PIXEL_SIZE && h_count < i_worm_x[17219:17214] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17219:17214] * PIXEL_SIZE && v_count < i_worm_y[17219:17214] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2870 < i_size && h_count >= i_worm_x[17225:17220] * PIXEL_SIZE && h_count < i_worm_x[17225:17220] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17225:17220] * PIXEL_SIZE && v_count < i_worm_y[17225:17220] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2871 < i_size && h_count >= i_worm_x[17231:17226] * PIXEL_SIZE && h_count < i_worm_x[17231:17226] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17231:17226] * PIXEL_SIZE && v_count < i_worm_y[17231:17226] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2872 < i_size && h_count >= i_worm_x[17237:17232] * PIXEL_SIZE && h_count < i_worm_x[17237:17232] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17237:17232] * PIXEL_SIZE && v_count < i_worm_y[17237:17232] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2873 < i_size && h_count >= i_worm_x[17243:17238] * PIXEL_SIZE && h_count < i_worm_x[17243:17238] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17243:17238] * PIXEL_SIZE && v_count < i_worm_y[17243:17238] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2874 < i_size && h_count >= i_worm_x[17249:17244] * PIXEL_SIZE && h_count < i_worm_x[17249:17244] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17249:17244] * PIXEL_SIZE && v_count < i_worm_y[17249:17244] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2875 < i_size && h_count >= i_worm_x[17255:17250] * PIXEL_SIZE && h_count < i_worm_x[17255:17250] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17255:17250] * PIXEL_SIZE && v_count < i_worm_y[17255:17250] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2876 < i_size && h_count >= i_worm_x[17261:17256] * PIXEL_SIZE && h_count < i_worm_x[17261:17256] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17261:17256] * PIXEL_SIZE && v_count < i_worm_y[17261:17256] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2877 < i_size && h_count >= i_worm_x[17267:17262] * PIXEL_SIZE && h_count < i_worm_x[17267:17262] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17267:17262] * PIXEL_SIZE && v_count < i_worm_y[17267:17262] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2878 < i_size && h_count >= i_worm_x[17273:17268] * PIXEL_SIZE && h_count < i_worm_x[17273:17268] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17273:17268] * PIXEL_SIZE && v_count < i_worm_y[17273:17268] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2879 < i_size && h_count >= i_worm_x[17279:17274] * PIXEL_SIZE && h_count < i_worm_x[17279:17274] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17279:17274] * PIXEL_SIZE && v_count < i_worm_y[17279:17274] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2880 < i_size && h_count >= i_worm_x[17285:17280] * PIXEL_SIZE && h_count < i_worm_x[17285:17280] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17285:17280] * PIXEL_SIZE && v_count < i_worm_y[17285:17280] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2881 < i_size && h_count >= i_worm_x[17291:17286] * PIXEL_SIZE && h_count < i_worm_x[17291:17286] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17291:17286] * PIXEL_SIZE && v_count < i_worm_y[17291:17286] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2882 < i_size && h_count >= i_worm_x[17297:17292] * PIXEL_SIZE && h_count < i_worm_x[17297:17292] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17297:17292] * PIXEL_SIZE && v_count < i_worm_y[17297:17292] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2883 < i_size && h_count >= i_worm_x[17303:17298] * PIXEL_SIZE && h_count < i_worm_x[17303:17298] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17303:17298] * PIXEL_SIZE && v_count < i_worm_y[17303:17298] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2884 < i_size && h_count >= i_worm_x[17309:17304] * PIXEL_SIZE && h_count < i_worm_x[17309:17304] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17309:17304] * PIXEL_SIZE && v_count < i_worm_y[17309:17304] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2885 < i_size && h_count >= i_worm_x[17315:17310] * PIXEL_SIZE && h_count < i_worm_x[17315:17310] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17315:17310] * PIXEL_SIZE && v_count < i_worm_y[17315:17310] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2886 < i_size && h_count >= i_worm_x[17321:17316] * PIXEL_SIZE && h_count < i_worm_x[17321:17316] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17321:17316] * PIXEL_SIZE && v_count < i_worm_y[17321:17316] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2887 < i_size && h_count >= i_worm_x[17327:17322] * PIXEL_SIZE && h_count < i_worm_x[17327:17322] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17327:17322] * PIXEL_SIZE && v_count < i_worm_y[17327:17322] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2888 < i_size && h_count >= i_worm_x[17333:17328] * PIXEL_SIZE && h_count < i_worm_x[17333:17328] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17333:17328] * PIXEL_SIZE && v_count < i_worm_y[17333:17328] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2889 < i_size && h_count >= i_worm_x[17339:17334] * PIXEL_SIZE && h_count < i_worm_x[17339:17334] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17339:17334] * PIXEL_SIZE && v_count < i_worm_y[17339:17334] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2890 < i_size && h_count >= i_worm_x[17345:17340] * PIXEL_SIZE && h_count < i_worm_x[17345:17340] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17345:17340] * PIXEL_SIZE && v_count < i_worm_y[17345:17340] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2891 < i_size && h_count >= i_worm_x[17351:17346] * PIXEL_SIZE && h_count < i_worm_x[17351:17346] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17351:17346] * PIXEL_SIZE && v_count < i_worm_y[17351:17346] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2892 < i_size && h_count >= i_worm_x[17357:17352] * PIXEL_SIZE && h_count < i_worm_x[17357:17352] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17357:17352] * PIXEL_SIZE && v_count < i_worm_y[17357:17352] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2893 < i_size && h_count >= i_worm_x[17363:17358] * PIXEL_SIZE && h_count < i_worm_x[17363:17358] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17363:17358] * PIXEL_SIZE && v_count < i_worm_y[17363:17358] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2894 < i_size && h_count >= i_worm_x[17369:17364] * PIXEL_SIZE && h_count < i_worm_x[17369:17364] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17369:17364] * PIXEL_SIZE && v_count < i_worm_y[17369:17364] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2895 < i_size && h_count >= i_worm_x[17375:17370] * PIXEL_SIZE && h_count < i_worm_x[17375:17370] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17375:17370] * PIXEL_SIZE && v_count < i_worm_y[17375:17370] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2896 < i_size && h_count >= i_worm_x[17381:17376] * PIXEL_SIZE && h_count < i_worm_x[17381:17376] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17381:17376] * PIXEL_SIZE && v_count < i_worm_y[17381:17376] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2897 < i_size && h_count >= i_worm_x[17387:17382] * PIXEL_SIZE && h_count < i_worm_x[17387:17382] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17387:17382] * PIXEL_SIZE && v_count < i_worm_y[17387:17382] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2898 < i_size && h_count >= i_worm_x[17393:17388] * PIXEL_SIZE && h_count < i_worm_x[17393:17388] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17393:17388] * PIXEL_SIZE && v_count < i_worm_y[17393:17388] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2899 < i_size && h_count >= i_worm_x[17399:17394] * PIXEL_SIZE && h_count < i_worm_x[17399:17394] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17399:17394] * PIXEL_SIZE && v_count < i_worm_y[17399:17394] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2900 < i_size && h_count >= i_worm_x[17405:17400] * PIXEL_SIZE && h_count < i_worm_x[17405:17400] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17405:17400] * PIXEL_SIZE && v_count < i_worm_y[17405:17400] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2901 < i_size && h_count >= i_worm_x[17411:17406] * PIXEL_SIZE && h_count < i_worm_x[17411:17406] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17411:17406] * PIXEL_SIZE && v_count < i_worm_y[17411:17406] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2902 < i_size && h_count >= i_worm_x[17417:17412] * PIXEL_SIZE && h_count < i_worm_x[17417:17412] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17417:17412] * PIXEL_SIZE && v_count < i_worm_y[17417:17412] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2903 < i_size && h_count >= i_worm_x[17423:17418] * PIXEL_SIZE && h_count < i_worm_x[17423:17418] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17423:17418] * PIXEL_SIZE && v_count < i_worm_y[17423:17418] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2904 < i_size && h_count >= i_worm_x[17429:17424] * PIXEL_SIZE && h_count < i_worm_x[17429:17424] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17429:17424] * PIXEL_SIZE && v_count < i_worm_y[17429:17424] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2905 < i_size && h_count >= i_worm_x[17435:17430] * PIXEL_SIZE && h_count < i_worm_x[17435:17430] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17435:17430] * PIXEL_SIZE && v_count < i_worm_y[17435:17430] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2906 < i_size && h_count >= i_worm_x[17441:17436] * PIXEL_SIZE && h_count < i_worm_x[17441:17436] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17441:17436] * PIXEL_SIZE && v_count < i_worm_y[17441:17436] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2907 < i_size && h_count >= i_worm_x[17447:17442] * PIXEL_SIZE && h_count < i_worm_x[17447:17442] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17447:17442] * PIXEL_SIZE && v_count < i_worm_y[17447:17442] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2908 < i_size && h_count >= i_worm_x[17453:17448] * PIXEL_SIZE && h_count < i_worm_x[17453:17448] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17453:17448] * PIXEL_SIZE && v_count < i_worm_y[17453:17448] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2909 < i_size && h_count >= i_worm_x[17459:17454] * PIXEL_SIZE && h_count < i_worm_x[17459:17454] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17459:17454] * PIXEL_SIZE && v_count < i_worm_y[17459:17454] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2910 < i_size && h_count >= i_worm_x[17465:17460] * PIXEL_SIZE && h_count < i_worm_x[17465:17460] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17465:17460] * PIXEL_SIZE && v_count < i_worm_y[17465:17460] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2911 < i_size && h_count >= i_worm_x[17471:17466] * PIXEL_SIZE && h_count < i_worm_x[17471:17466] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17471:17466] * PIXEL_SIZE && v_count < i_worm_y[17471:17466] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2912 < i_size && h_count >= i_worm_x[17477:17472] * PIXEL_SIZE && h_count < i_worm_x[17477:17472] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17477:17472] * PIXEL_SIZE && v_count < i_worm_y[17477:17472] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2913 < i_size && h_count >= i_worm_x[17483:17478] * PIXEL_SIZE && h_count < i_worm_x[17483:17478] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17483:17478] * PIXEL_SIZE && v_count < i_worm_y[17483:17478] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2914 < i_size && h_count >= i_worm_x[17489:17484] * PIXEL_SIZE && h_count < i_worm_x[17489:17484] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17489:17484] * PIXEL_SIZE && v_count < i_worm_y[17489:17484] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2915 < i_size && h_count >= i_worm_x[17495:17490] * PIXEL_SIZE && h_count < i_worm_x[17495:17490] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17495:17490] * PIXEL_SIZE && v_count < i_worm_y[17495:17490] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2916 < i_size && h_count >= i_worm_x[17501:17496] * PIXEL_SIZE && h_count < i_worm_x[17501:17496] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17501:17496] * PIXEL_SIZE && v_count < i_worm_y[17501:17496] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2917 < i_size && h_count >= i_worm_x[17507:17502] * PIXEL_SIZE && h_count < i_worm_x[17507:17502] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17507:17502] * PIXEL_SIZE && v_count < i_worm_y[17507:17502] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2918 < i_size && h_count >= i_worm_x[17513:17508] * PIXEL_SIZE && h_count < i_worm_x[17513:17508] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17513:17508] * PIXEL_SIZE && v_count < i_worm_y[17513:17508] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2919 < i_size && h_count >= i_worm_x[17519:17514] * PIXEL_SIZE && h_count < i_worm_x[17519:17514] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17519:17514] * PIXEL_SIZE && v_count < i_worm_y[17519:17514] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2920 < i_size && h_count >= i_worm_x[17525:17520] * PIXEL_SIZE && h_count < i_worm_x[17525:17520] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17525:17520] * PIXEL_SIZE && v_count < i_worm_y[17525:17520] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2921 < i_size && h_count >= i_worm_x[17531:17526] * PIXEL_SIZE && h_count < i_worm_x[17531:17526] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17531:17526] * PIXEL_SIZE && v_count < i_worm_y[17531:17526] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2922 < i_size && h_count >= i_worm_x[17537:17532] * PIXEL_SIZE && h_count < i_worm_x[17537:17532] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17537:17532] * PIXEL_SIZE && v_count < i_worm_y[17537:17532] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2923 < i_size && h_count >= i_worm_x[17543:17538] * PIXEL_SIZE && h_count < i_worm_x[17543:17538] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17543:17538] * PIXEL_SIZE && v_count < i_worm_y[17543:17538] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2924 < i_size && h_count >= i_worm_x[17549:17544] * PIXEL_SIZE && h_count < i_worm_x[17549:17544] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17549:17544] * PIXEL_SIZE && v_count < i_worm_y[17549:17544] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2925 < i_size && h_count >= i_worm_x[17555:17550] * PIXEL_SIZE && h_count < i_worm_x[17555:17550] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17555:17550] * PIXEL_SIZE && v_count < i_worm_y[17555:17550] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2926 < i_size && h_count >= i_worm_x[17561:17556] * PIXEL_SIZE && h_count < i_worm_x[17561:17556] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17561:17556] * PIXEL_SIZE && v_count < i_worm_y[17561:17556] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2927 < i_size && h_count >= i_worm_x[17567:17562] * PIXEL_SIZE && h_count < i_worm_x[17567:17562] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17567:17562] * PIXEL_SIZE && v_count < i_worm_y[17567:17562] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2928 < i_size && h_count >= i_worm_x[17573:17568] * PIXEL_SIZE && h_count < i_worm_x[17573:17568] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17573:17568] * PIXEL_SIZE && v_count < i_worm_y[17573:17568] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2929 < i_size && h_count >= i_worm_x[17579:17574] * PIXEL_SIZE && h_count < i_worm_x[17579:17574] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17579:17574] * PIXEL_SIZE && v_count < i_worm_y[17579:17574] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2930 < i_size && h_count >= i_worm_x[17585:17580] * PIXEL_SIZE && h_count < i_worm_x[17585:17580] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17585:17580] * PIXEL_SIZE && v_count < i_worm_y[17585:17580] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2931 < i_size && h_count >= i_worm_x[17591:17586] * PIXEL_SIZE && h_count < i_worm_x[17591:17586] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17591:17586] * PIXEL_SIZE && v_count < i_worm_y[17591:17586] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2932 < i_size && h_count >= i_worm_x[17597:17592] * PIXEL_SIZE && h_count < i_worm_x[17597:17592] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17597:17592] * PIXEL_SIZE && v_count < i_worm_y[17597:17592] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2933 < i_size && h_count >= i_worm_x[17603:17598] * PIXEL_SIZE && h_count < i_worm_x[17603:17598] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17603:17598] * PIXEL_SIZE && v_count < i_worm_y[17603:17598] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2934 < i_size && h_count >= i_worm_x[17609:17604] * PIXEL_SIZE && h_count < i_worm_x[17609:17604] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17609:17604] * PIXEL_SIZE && v_count < i_worm_y[17609:17604] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2935 < i_size && h_count >= i_worm_x[17615:17610] * PIXEL_SIZE && h_count < i_worm_x[17615:17610] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17615:17610] * PIXEL_SIZE && v_count < i_worm_y[17615:17610] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2936 < i_size && h_count >= i_worm_x[17621:17616] * PIXEL_SIZE && h_count < i_worm_x[17621:17616] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17621:17616] * PIXEL_SIZE && v_count < i_worm_y[17621:17616] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2937 < i_size && h_count >= i_worm_x[17627:17622] * PIXEL_SIZE && h_count < i_worm_x[17627:17622] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17627:17622] * PIXEL_SIZE && v_count < i_worm_y[17627:17622] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2938 < i_size && h_count >= i_worm_x[17633:17628] * PIXEL_SIZE && h_count < i_worm_x[17633:17628] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17633:17628] * PIXEL_SIZE && v_count < i_worm_y[17633:17628] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2939 < i_size && h_count >= i_worm_x[17639:17634] * PIXEL_SIZE && h_count < i_worm_x[17639:17634] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17639:17634] * PIXEL_SIZE && v_count < i_worm_y[17639:17634] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2940 < i_size && h_count >= i_worm_x[17645:17640] * PIXEL_SIZE && h_count < i_worm_x[17645:17640] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17645:17640] * PIXEL_SIZE && v_count < i_worm_y[17645:17640] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2941 < i_size && h_count >= i_worm_x[17651:17646] * PIXEL_SIZE && h_count < i_worm_x[17651:17646] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17651:17646] * PIXEL_SIZE && v_count < i_worm_y[17651:17646] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2942 < i_size && h_count >= i_worm_x[17657:17652] * PIXEL_SIZE && h_count < i_worm_x[17657:17652] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17657:17652] * PIXEL_SIZE && v_count < i_worm_y[17657:17652] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2943 < i_size && h_count >= i_worm_x[17663:17658] * PIXEL_SIZE && h_count < i_worm_x[17663:17658] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17663:17658] * PIXEL_SIZE && v_count < i_worm_y[17663:17658] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2944 < i_size && h_count >= i_worm_x[17669:17664] * PIXEL_SIZE && h_count < i_worm_x[17669:17664] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17669:17664] * PIXEL_SIZE && v_count < i_worm_y[17669:17664] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2945 < i_size && h_count >= i_worm_x[17675:17670] * PIXEL_SIZE && h_count < i_worm_x[17675:17670] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17675:17670] * PIXEL_SIZE && v_count < i_worm_y[17675:17670] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2946 < i_size && h_count >= i_worm_x[17681:17676] * PIXEL_SIZE && h_count < i_worm_x[17681:17676] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17681:17676] * PIXEL_SIZE && v_count < i_worm_y[17681:17676] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2947 < i_size && h_count >= i_worm_x[17687:17682] * PIXEL_SIZE && h_count < i_worm_x[17687:17682] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17687:17682] * PIXEL_SIZE && v_count < i_worm_y[17687:17682] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2948 < i_size && h_count >= i_worm_x[17693:17688] * PIXEL_SIZE && h_count < i_worm_x[17693:17688] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17693:17688] * PIXEL_SIZE && v_count < i_worm_y[17693:17688] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2949 < i_size && h_count >= i_worm_x[17699:17694] * PIXEL_SIZE && h_count < i_worm_x[17699:17694] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17699:17694] * PIXEL_SIZE && v_count < i_worm_y[17699:17694] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2950 < i_size && h_count >= i_worm_x[17705:17700] * PIXEL_SIZE && h_count < i_worm_x[17705:17700] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17705:17700] * PIXEL_SIZE && v_count < i_worm_y[17705:17700] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2951 < i_size && h_count >= i_worm_x[17711:17706] * PIXEL_SIZE && h_count < i_worm_x[17711:17706] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17711:17706] * PIXEL_SIZE && v_count < i_worm_y[17711:17706] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2952 < i_size && h_count >= i_worm_x[17717:17712] * PIXEL_SIZE && h_count < i_worm_x[17717:17712] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17717:17712] * PIXEL_SIZE && v_count < i_worm_y[17717:17712] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2953 < i_size && h_count >= i_worm_x[17723:17718] * PIXEL_SIZE && h_count < i_worm_x[17723:17718] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17723:17718] * PIXEL_SIZE && v_count < i_worm_y[17723:17718] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2954 < i_size && h_count >= i_worm_x[17729:17724] * PIXEL_SIZE && h_count < i_worm_x[17729:17724] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17729:17724] * PIXEL_SIZE && v_count < i_worm_y[17729:17724] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2955 < i_size && h_count >= i_worm_x[17735:17730] * PIXEL_SIZE && h_count < i_worm_x[17735:17730] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17735:17730] * PIXEL_SIZE && v_count < i_worm_y[17735:17730] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2956 < i_size && h_count >= i_worm_x[17741:17736] * PIXEL_SIZE && h_count < i_worm_x[17741:17736] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17741:17736] * PIXEL_SIZE && v_count < i_worm_y[17741:17736] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2957 < i_size && h_count >= i_worm_x[17747:17742] * PIXEL_SIZE && h_count < i_worm_x[17747:17742] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17747:17742] * PIXEL_SIZE && v_count < i_worm_y[17747:17742] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2958 < i_size && h_count >= i_worm_x[17753:17748] * PIXEL_SIZE && h_count < i_worm_x[17753:17748] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17753:17748] * PIXEL_SIZE && v_count < i_worm_y[17753:17748] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2959 < i_size && h_count >= i_worm_x[17759:17754] * PIXEL_SIZE && h_count < i_worm_x[17759:17754] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17759:17754] * PIXEL_SIZE && v_count < i_worm_y[17759:17754] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2960 < i_size && h_count >= i_worm_x[17765:17760] * PIXEL_SIZE && h_count < i_worm_x[17765:17760] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17765:17760] * PIXEL_SIZE && v_count < i_worm_y[17765:17760] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2961 < i_size && h_count >= i_worm_x[17771:17766] * PIXEL_SIZE && h_count < i_worm_x[17771:17766] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17771:17766] * PIXEL_SIZE && v_count < i_worm_y[17771:17766] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2962 < i_size && h_count >= i_worm_x[17777:17772] * PIXEL_SIZE && h_count < i_worm_x[17777:17772] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17777:17772] * PIXEL_SIZE && v_count < i_worm_y[17777:17772] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2963 < i_size && h_count >= i_worm_x[17783:17778] * PIXEL_SIZE && h_count < i_worm_x[17783:17778] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17783:17778] * PIXEL_SIZE && v_count < i_worm_y[17783:17778] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2964 < i_size && h_count >= i_worm_x[17789:17784] * PIXEL_SIZE && h_count < i_worm_x[17789:17784] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17789:17784] * PIXEL_SIZE && v_count < i_worm_y[17789:17784] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2965 < i_size && h_count >= i_worm_x[17795:17790] * PIXEL_SIZE && h_count < i_worm_x[17795:17790] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17795:17790] * PIXEL_SIZE && v_count < i_worm_y[17795:17790] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2966 < i_size && h_count >= i_worm_x[17801:17796] * PIXEL_SIZE && h_count < i_worm_x[17801:17796] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17801:17796] * PIXEL_SIZE && v_count < i_worm_y[17801:17796] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2967 < i_size && h_count >= i_worm_x[17807:17802] * PIXEL_SIZE && h_count < i_worm_x[17807:17802] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17807:17802] * PIXEL_SIZE && v_count < i_worm_y[17807:17802] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2968 < i_size && h_count >= i_worm_x[17813:17808] * PIXEL_SIZE && h_count < i_worm_x[17813:17808] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17813:17808] * PIXEL_SIZE && v_count < i_worm_y[17813:17808] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2969 < i_size && h_count >= i_worm_x[17819:17814] * PIXEL_SIZE && h_count < i_worm_x[17819:17814] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17819:17814] * PIXEL_SIZE && v_count < i_worm_y[17819:17814] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2970 < i_size && h_count >= i_worm_x[17825:17820] * PIXEL_SIZE && h_count < i_worm_x[17825:17820] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17825:17820] * PIXEL_SIZE && v_count < i_worm_y[17825:17820] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2971 < i_size && h_count >= i_worm_x[17831:17826] * PIXEL_SIZE && h_count < i_worm_x[17831:17826] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17831:17826] * PIXEL_SIZE && v_count < i_worm_y[17831:17826] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2972 < i_size && h_count >= i_worm_x[17837:17832] * PIXEL_SIZE && h_count < i_worm_x[17837:17832] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17837:17832] * PIXEL_SIZE && v_count < i_worm_y[17837:17832] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2973 < i_size && h_count >= i_worm_x[17843:17838] * PIXEL_SIZE && h_count < i_worm_x[17843:17838] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17843:17838] * PIXEL_SIZE && v_count < i_worm_y[17843:17838] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2974 < i_size && h_count >= i_worm_x[17849:17844] * PIXEL_SIZE && h_count < i_worm_x[17849:17844] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17849:17844] * PIXEL_SIZE && v_count < i_worm_y[17849:17844] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2975 < i_size && h_count >= i_worm_x[17855:17850] * PIXEL_SIZE && h_count < i_worm_x[17855:17850] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17855:17850] * PIXEL_SIZE && v_count < i_worm_y[17855:17850] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2976 < i_size && h_count >= i_worm_x[17861:17856] * PIXEL_SIZE && h_count < i_worm_x[17861:17856] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17861:17856] * PIXEL_SIZE && v_count < i_worm_y[17861:17856] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2977 < i_size && h_count >= i_worm_x[17867:17862] * PIXEL_SIZE && h_count < i_worm_x[17867:17862] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17867:17862] * PIXEL_SIZE && v_count < i_worm_y[17867:17862] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2978 < i_size && h_count >= i_worm_x[17873:17868] * PIXEL_SIZE && h_count < i_worm_x[17873:17868] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17873:17868] * PIXEL_SIZE && v_count < i_worm_y[17873:17868] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2979 < i_size && h_count >= i_worm_x[17879:17874] * PIXEL_SIZE && h_count < i_worm_x[17879:17874] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17879:17874] * PIXEL_SIZE && v_count < i_worm_y[17879:17874] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2980 < i_size && h_count >= i_worm_x[17885:17880] * PIXEL_SIZE && h_count < i_worm_x[17885:17880] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17885:17880] * PIXEL_SIZE && v_count < i_worm_y[17885:17880] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2981 < i_size && h_count >= i_worm_x[17891:17886] * PIXEL_SIZE && h_count < i_worm_x[17891:17886] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17891:17886] * PIXEL_SIZE && v_count < i_worm_y[17891:17886] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2982 < i_size && h_count >= i_worm_x[17897:17892] * PIXEL_SIZE && h_count < i_worm_x[17897:17892] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17897:17892] * PIXEL_SIZE && v_count < i_worm_y[17897:17892] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2983 < i_size && h_count >= i_worm_x[17903:17898] * PIXEL_SIZE && h_count < i_worm_x[17903:17898] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17903:17898] * PIXEL_SIZE && v_count < i_worm_y[17903:17898] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2984 < i_size && h_count >= i_worm_x[17909:17904] * PIXEL_SIZE && h_count < i_worm_x[17909:17904] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17909:17904] * PIXEL_SIZE && v_count < i_worm_y[17909:17904] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2985 < i_size && h_count >= i_worm_x[17915:17910] * PIXEL_SIZE && h_count < i_worm_x[17915:17910] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17915:17910] * PIXEL_SIZE && v_count < i_worm_y[17915:17910] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2986 < i_size && h_count >= i_worm_x[17921:17916] * PIXEL_SIZE && h_count < i_worm_x[17921:17916] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17921:17916] * PIXEL_SIZE && v_count < i_worm_y[17921:17916] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2987 < i_size && h_count >= i_worm_x[17927:17922] * PIXEL_SIZE && h_count < i_worm_x[17927:17922] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17927:17922] * PIXEL_SIZE && v_count < i_worm_y[17927:17922] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2988 < i_size && h_count >= i_worm_x[17933:17928] * PIXEL_SIZE && h_count < i_worm_x[17933:17928] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17933:17928] * PIXEL_SIZE && v_count < i_worm_y[17933:17928] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2989 < i_size && h_count >= i_worm_x[17939:17934] * PIXEL_SIZE && h_count < i_worm_x[17939:17934] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17939:17934] * PIXEL_SIZE && v_count < i_worm_y[17939:17934] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2990 < i_size && h_count >= i_worm_x[17945:17940] * PIXEL_SIZE && h_count < i_worm_x[17945:17940] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17945:17940] * PIXEL_SIZE && v_count < i_worm_y[17945:17940] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2991 < i_size && h_count >= i_worm_x[17951:17946] * PIXEL_SIZE && h_count < i_worm_x[17951:17946] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17951:17946] * PIXEL_SIZE && v_count < i_worm_y[17951:17946] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2992 < i_size && h_count >= i_worm_x[17957:17952] * PIXEL_SIZE && h_count < i_worm_x[17957:17952] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17957:17952] * PIXEL_SIZE && v_count < i_worm_y[17957:17952] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2993 < i_size && h_count >= i_worm_x[17963:17958] * PIXEL_SIZE && h_count < i_worm_x[17963:17958] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17963:17958] * PIXEL_SIZE && v_count < i_worm_y[17963:17958] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2994 < i_size && h_count >= i_worm_x[17969:17964] * PIXEL_SIZE && h_count < i_worm_x[17969:17964] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17969:17964] * PIXEL_SIZE && v_count < i_worm_y[17969:17964] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2995 < i_size && h_count >= i_worm_x[17975:17970] * PIXEL_SIZE && h_count < i_worm_x[17975:17970] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17975:17970] * PIXEL_SIZE && v_count < i_worm_y[17975:17970] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2996 < i_size && h_count >= i_worm_x[17981:17976] * PIXEL_SIZE && h_count < i_worm_x[17981:17976] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17981:17976] * PIXEL_SIZE && v_count < i_worm_y[17981:17976] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2997 < i_size && h_count >= i_worm_x[17987:17982] * PIXEL_SIZE && h_count < i_worm_x[17987:17982] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17987:17982] * PIXEL_SIZE && v_count < i_worm_y[17987:17982] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2998 < i_size && h_count >= i_worm_x[17993:17988] * PIXEL_SIZE && h_count < i_worm_x[17993:17988] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17993:17988] * PIXEL_SIZE && v_count < i_worm_y[17993:17988] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (2999 < i_size && h_count >= i_worm_x[17999:17994] * PIXEL_SIZE && h_count < i_worm_x[17999:17994] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[17999:17994] * PIXEL_SIZE && v_count < i_worm_y[17999:17994] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3000 < i_size && h_count >= i_worm_x[18005:18000] * PIXEL_SIZE && h_count < i_worm_x[18005:18000] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18005:18000] * PIXEL_SIZE && v_count < i_worm_y[18005:18000] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3001 < i_size && h_count >= i_worm_x[18011:18006] * PIXEL_SIZE && h_count < i_worm_x[18011:18006] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18011:18006] * PIXEL_SIZE && v_count < i_worm_y[18011:18006] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3002 < i_size && h_count >= i_worm_x[18017:18012] * PIXEL_SIZE && h_count < i_worm_x[18017:18012] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18017:18012] * PIXEL_SIZE && v_count < i_worm_y[18017:18012] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3003 < i_size && h_count >= i_worm_x[18023:18018] * PIXEL_SIZE && h_count < i_worm_x[18023:18018] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18023:18018] * PIXEL_SIZE && v_count < i_worm_y[18023:18018] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3004 < i_size && h_count >= i_worm_x[18029:18024] * PIXEL_SIZE && h_count < i_worm_x[18029:18024] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18029:18024] * PIXEL_SIZE && v_count < i_worm_y[18029:18024] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3005 < i_size && h_count >= i_worm_x[18035:18030] * PIXEL_SIZE && h_count < i_worm_x[18035:18030] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18035:18030] * PIXEL_SIZE && v_count < i_worm_y[18035:18030] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3006 < i_size && h_count >= i_worm_x[18041:18036] * PIXEL_SIZE && h_count < i_worm_x[18041:18036] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18041:18036] * PIXEL_SIZE && v_count < i_worm_y[18041:18036] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3007 < i_size && h_count >= i_worm_x[18047:18042] * PIXEL_SIZE && h_count < i_worm_x[18047:18042] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18047:18042] * PIXEL_SIZE && v_count < i_worm_y[18047:18042] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3008 < i_size && h_count >= i_worm_x[18053:18048] * PIXEL_SIZE && h_count < i_worm_x[18053:18048] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18053:18048] * PIXEL_SIZE && v_count < i_worm_y[18053:18048] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3009 < i_size && h_count >= i_worm_x[18059:18054] * PIXEL_SIZE && h_count < i_worm_x[18059:18054] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18059:18054] * PIXEL_SIZE && v_count < i_worm_y[18059:18054] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3010 < i_size && h_count >= i_worm_x[18065:18060] * PIXEL_SIZE && h_count < i_worm_x[18065:18060] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18065:18060] * PIXEL_SIZE && v_count < i_worm_y[18065:18060] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3011 < i_size && h_count >= i_worm_x[18071:18066] * PIXEL_SIZE && h_count < i_worm_x[18071:18066] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18071:18066] * PIXEL_SIZE && v_count < i_worm_y[18071:18066] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3012 < i_size && h_count >= i_worm_x[18077:18072] * PIXEL_SIZE && h_count < i_worm_x[18077:18072] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18077:18072] * PIXEL_SIZE && v_count < i_worm_y[18077:18072] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3013 < i_size && h_count >= i_worm_x[18083:18078] * PIXEL_SIZE && h_count < i_worm_x[18083:18078] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18083:18078] * PIXEL_SIZE && v_count < i_worm_y[18083:18078] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3014 < i_size && h_count >= i_worm_x[18089:18084] * PIXEL_SIZE && h_count < i_worm_x[18089:18084] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18089:18084] * PIXEL_SIZE && v_count < i_worm_y[18089:18084] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3015 < i_size && h_count >= i_worm_x[18095:18090] * PIXEL_SIZE && h_count < i_worm_x[18095:18090] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18095:18090] * PIXEL_SIZE && v_count < i_worm_y[18095:18090] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3016 < i_size && h_count >= i_worm_x[18101:18096] * PIXEL_SIZE && h_count < i_worm_x[18101:18096] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18101:18096] * PIXEL_SIZE && v_count < i_worm_y[18101:18096] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3017 < i_size && h_count >= i_worm_x[18107:18102] * PIXEL_SIZE && h_count < i_worm_x[18107:18102] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18107:18102] * PIXEL_SIZE && v_count < i_worm_y[18107:18102] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3018 < i_size && h_count >= i_worm_x[18113:18108] * PIXEL_SIZE && h_count < i_worm_x[18113:18108] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18113:18108] * PIXEL_SIZE && v_count < i_worm_y[18113:18108] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3019 < i_size && h_count >= i_worm_x[18119:18114] * PIXEL_SIZE && h_count < i_worm_x[18119:18114] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18119:18114] * PIXEL_SIZE && v_count < i_worm_y[18119:18114] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3020 < i_size && h_count >= i_worm_x[18125:18120] * PIXEL_SIZE && h_count < i_worm_x[18125:18120] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18125:18120] * PIXEL_SIZE && v_count < i_worm_y[18125:18120] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3021 < i_size && h_count >= i_worm_x[18131:18126] * PIXEL_SIZE && h_count < i_worm_x[18131:18126] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18131:18126] * PIXEL_SIZE && v_count < i_worm_y[18131:18126] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3022 < i_size && h_count >= i_worm_x[18137:18132] * PIXEL_SIZE && h_count < i_worm_x[18137:18132] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18137:18132] * PIXEL_SIZE && v_count < i_worm_y[18137:18132] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3023 < i_size && h_count >= i_worm_x[18143:18138] * PIXEL_SIZE && h_count < i_worm_x[18143:18138] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18143:18138] * PIXEL_SIZE && v_count < i_worm_y[18143:18138] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3024 < i_size && h_count >= i_worm_x[18149:18144] * PIXEL_SIZE && h_count < i_worm_x[18149:18144] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18149:18144] * PIXEL_SIZE && v_count < i_worm_y[18149:18144] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3025 < i_size && h_count >= i_worm_x[18155:18150] * PIXEL_SIZE && h_count < i_worm_x[18155:18150] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18155:18150] * PIXEL_SIZE && v_count < i_worm_y[18155:18150] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3026 < i_size && h_count >= i_worm_x[18161:18156] * PIXEL_SIZE && h_count < i_worm_x[18161:18156] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18161:18156] * PIXEL_SIZE && v_count < i_worm_y[18161:18156] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3027 < i_size && h_count >= i_worm_x[18167:18162] * PIXEL_SIZE && h_count < i_worm_x[18167:18162] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18167:18162] * PIXEL_SIZE && v_count < i_worm_y[18167:18162] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3028 < i_size && h_count >= i_worm_x[18173:18168] * PIXEL_SIZE && h_count < i_worm_x[18173:18168] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18173:18168] * PIXEL_SIZE && v_count < i_worm_y[18173:18168] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3029 < i_size && h_count >= i_worm_x[18179:18174] * PIXEL_SIZE && h_count < i_worm_x[18179:18174] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18179:18174] * PIXEL_SIZE && v_count < i_worm_y[18179:18174] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3030 < i_size && h_count >= i_worm_x[18185:18180] * PIXEL_SIZE && h_count < i_worm_x[18185:18180] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18185:18180] * PIXEL_SIZE && v_count < i_worm_y[18185:18180] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3031 < i_size && h_count >= i_worm_x[18191:18186] * PIXEL_SIZE && h_count < i_worm_x[18191:18186] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18191:18186] * PIXEL_SIZE && v_count < i_worm_y[18191:18186] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3032 < i_size && h_count >= i_worm_x[18197:18192] * PIXEL_SIZE && h_count < i_worm_x[18197:18192] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18197:18192] * PIXEL_SIZE && v_count < i_worm_y[18197:18192] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3033 < i_size && h_count >= i_worm_x[18203:18198] * PIXEL_SIZE && h_count < i_worm_x[18203:18198] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18203:18198] * PIXEL_SIZE && v_count < i_worm_y[18203:18198] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3034 < i_size && h_count >= i_worm_x[18209:18204] * PIXEL_SIZE && h_count < i_worm_x[18209:18204] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18209:18204] * PIXEL_SIZE && v_count < i_worm_y[18209:18204] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3035 < i_size && h_count >= i_worm_x[18215:18210] * PIXEL_SIZE && h_count < i_worm_x[18215:18210] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18215:18210] * PIXEL_SIZE && v_count < i_worm_y[18215:18210] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3036 < i_size && h_count >= i_worm_x[18221:18216] * PIXEL_SIZE && h_count < i_worm_x[18221:18216] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18221:18216] * PIXEL_SIZE && v_count < i_worm_y[18221:18216] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3037 < i_size && h_count >= i_worm_x[18227:18222] * PIXEL_SIZE && h_count < i_worm_x[18227:18222] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18227:18222] * PIXEL_SIZE && v_count < i_worm_y[18227:18222] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3038 < i_size && h_count >= i_worm_x[18233:18228] * PIXEL_SIZE && h_count < i_worm_x[18233:18228] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18233:18228] * PIXEL_SIZE && v_count < i_worm_y[18233:18228] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3039 < i_size && h_count >= i_worm_x[18239:18234] * PIXEL_SIZE && h_count < i_worm_x[18239:18234] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18239:18234] * PIXEL_SIZE && v_count < i_worm_y[18239:18234] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3040 < i_size && h_count >= i_worm_x[18245:18240] * PIXEL_SIZE && h_count < i_worm_x[18245:18240] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18245:18240] * PIXEL_SIZE && v_count < i_worm_y[18245:18240] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3041 < i_size && h_count >= i_worm_x[18251:18246] * PIXEL_SIZE && h_count < i_worm_x[18251:18246] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18251:18246] * PIXEL_SIZE && v_count < i_worm_y[18251:18246] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3042 < i_size && h_count >= i_worm_x[18257:18252] * PIXEL_SIZE && h_count < i_worm_x[18257:18252] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18257:18252] * PIXEL_SIZE && v_count < i_worm_y[18257:18252] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3043 < i_size && h_count >= i_worm_x[18263:18258] * PIXEL_SIZE && h_count < i_worm_x[18263:18258] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18263:18258] * PIXEL_SIZE && v_count < i_worm_y[18263:18258] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3044 < i_size && h_count >= i_worm_x[18269:18264] * PIXEL_SIZE && h_count < i_worm_x[18269:18264] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18269:18264] * PIXEL_SIZE && v_count < i_worm_y[18269:18264] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3045 < i_size && h_count >= i_worm_x[18275:18270] * PIXEL_SIZE && h_count < i_worm_x[18275:18270] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18275:18270] * PIXEL_SIZE && v_count < i_worm_y[18275:18270] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3046 < i_size && h_count >= i_worm_x[18281:18276] * PIXEL_SIZE && h_count < i_worm_x[18281:18276] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18281:18276] * PIXEL_SIZE && v_count < i_worm_y[18281:18276] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3047 < i_size && h_count >= i_worm_x[18287:18282] * PIXEL_SIZE && h_count < i_worm_x[18287:18282] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18287:18282] * PIXEL_SIZE && v_count < i_worm_y[18287:18282] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3048 < i_size && h_count >= i_worm_x[18293:18288] * PIXEL_SIZE && h_count < i_worm_x[18293:18288] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18293:18288] * PIXEL_SIZE && v_count < i_worm_y[18293:18288] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3049 < i_size && h_count >= i_worm_x[18299:18294] * PIXEL_SIZE && h_count < i_worm_x[18299:18294] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18299:18294] * PIXEL_SIZE && v_count < i_worm_y[18299:18294] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3050 < i_size && h_count >= i_worm_x[18305:18300] * PIXEL_SIZE && h_count < i_worm_x[18305:18300] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18305:18300] * PIXEL_SIZE && v_count < i_worm_y[18305:18300] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3051 < i_size && h_count >= i_worm_x[18311:18306] * PIXEL_SIZE && h_count < i_worm_x[18311:18306] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18311:18306] * PIXEL_SIZE && v_count < i_worm_y[18311:18306] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3052 < i_size && h_count >= i_worm_x[18317:18312] * PIXEL_SIZE && h_count < i_worm_x[18317:18312] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18317:18312] * PIXEL_SIZE && v_count < i_worm_y[18317:18312] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3053 < i_size && h_count >= i_worm_x[18323:18318] * PIXEL_SIZE && h_count < i_worm_x[18323:18318] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18323:18318] * PIXEL_SIZE && v_count < i_worm_y[18323:18318] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3054 < i_size && h_count >= i_worm_x[18329:18324] * PIXEL_SIZE && h_count < i_worm_x[18329:18324] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18329:18324] * PIXEL_SIZE && v_count < i_worm_y[18329:18324] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3055 < i_size && h_count >= i_worm_x[18335:18330] * PIXEL_SIZE && h_count < i_worm_x[18335:18330] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18335:18330] * PIXEL_SIZE && v_count < i_worm_y[18335:18330] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3056 < i_size && h_count >= i_worm_x[18341:18336] * PIXEL_SIZE && h_count < i_worm_x[18341:18336] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18341:18336] * PIXEL_SIZE && v_count < i_worm_y[18341:18336] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3057 < i_size && h_count >= i_worm_x[18347:18342] * PIXEL_SIZE && h_count < i_worm_x[18347:18342] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18347:18342] * PIXEL_SIZE && v_count < i_worm_y[18347:18342] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3058 < i_size && h_count >= i_worm_x[18353:18348] * PIXEL_SIZE && h_count < i_worm_x[18353:18348] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18353:18348] * PIXEL_SIZE && v_count < i_worm_y[18353:18348] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3059 < i_size && h_count >= i_worm_x[18359:18354] * PIXEL_SIZE && h_count < i_worm_x[18359:18354] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18359:18354] * PIXEL_SIZE && v_count < i_worm_y[18359:18354] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3060 < i_size && h_count >= i_worm_x[18365:18360] * PIXEL_SIZE && h_count < i_worm_x[18365:18360] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18365:18360] * PIXEL_SIZE && v_count < i_worm_y[18365:18360] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3061 < i_size && h_count >= i_worm_x[18371:18366] * PIXEL_SIZE && h_count < i_worm_x[18371:18366] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18371:18366] * PIXEL_SIZE && v_count < i_worm_y[18371:18366] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3062 < i_size && h_count >= i_worm_x[18377:18372] * PIXEL_SIZE && h_count < i_worm_x[18377:18372] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18377:18372] * PIXEL_SIZE && v_count < i_worm_y[18377:18372] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3063 < i_size && h_count >= i_worm_x[18383:18378] * PIXEL_SIZE && h_count < i_worm_x[18383:18378] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18383:18378] * PIXEL_SIZE && v_count < i_worm_y[18383:18378] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3064 < i_size && h_count >= i_worm_x[18389:18384] * PIXEL_SIZE && h_count < i_worm_x[18389:18384] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18389:18384] * PIXEL_SIZE && v_count < i_worm_y[18389:18384] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3065 < i_size && h_count >= i_worm_x[18395:18390] * PIXEL_SIZE && h_count < i_worm_x[18395:18390] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18395:18390] * PIXEL_SIZE && v_count < i_worm_y[18395:18390] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3066 < i_size && h_count >= i_worm_x[18401:18396] * PIXEL_SIZE && h_count < i_worm_x[18401:18396] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18401:18396] * PIXEL_SIZE && v_count < i_worm_y[18401:18396] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3067 < i_size && h_count >= i_worm_x[18407:18402] * PIXEL_SIZE && h_count < i_worm_x[18407:18402] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18407:18402] * PIXEL_SIZE && v_count < i_worm_y[18407:18402] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3068 < i_size && h_count >= i_worm_x[18413:18408] * PIXEL_SIZE && h_count < i_worm_x[18413:18408] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18413:18408] * PIXEL_SIZE && v_count < i_worm_y[18413:18408] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3069 < i_size && h_count >= i_worm_x[18419:18414] * PIXEL_SIZE && h_count < i_worm_x[18419:18414] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18419:18414] * PIXEL_SIZE && v_count < i_worm_y[18419:18414] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3070 < i_size && h_count >= i_worm_x[18425:18420] * PIXEL_SIZE && h_count < i_worm_x[18425:18420] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18425:18420] * PIXEL_SIZE && v_count < i_worm_y[18425:18420] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end
                     if (3071 < i_size && h_count >= i_worm_x[18431:18426] * PIXEL_SIZE && h_count < i_worm_x[18431:18426] * PIXEL_SIZE + PIXEL_SIZE &&
                          v_count >= i_worm_y[18431:18426] * PIXEL_SIZE && v_count < i_worm_y[18431:18426] * PIXEL_SIZE + PIXEL_SIZE) begin
                      worm_active = 1;
                    end


                if (worm_active) begin
                    // 지렁이 위치 (빨강색)
                    o_red <= 8'hF;
                    o_green <= 8'h0;
                    o_blue <= 8'h0;
                end else if (item_active) begin
                    // 아이템 위치 (초록색)
                    o_red <= 8'h0;
                    o_green <= 8'hF;
                    o_blue <= 8'h0;
                end else if (edge_active) begin
                    // 가장자리 (흰색)
                    o_red <= 8'hF;
                    o_green <= 8'hF;
                    o_blue <= 8'hF;
                end else begin
                    // 나머지 영역 (검정색)
                    o_red <= 8'h0;
                    o_green <= 8'h0;
                    o_blue <= 8'h0;
                end
            end else begin
                // 640 * 480 영역 밖
                o_red <= 8'h0;
                o_green <= 8'h0;
                o_blue <= 8'h0;
            end
        end
    end
endmodule